VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sb_0__0_
  CLASS BLOCK ;
  FOREIGN sb_0__0_ ;
  ORIGIN 0.000 0.000 ;
  SIZE 100.000 BY 100.000 ;
  PIN ccff_head
    PORT
      LAYER met3 ;
        RECT 0.000 74.840 4.000 75.440 ;
    END
  END ccff_head
  PIN ccff_tail
    PORT
      LAYER met3 ;
        RECT 96.000 6.840 100.000 7.440 ;
    END
  END ccff_tail
  PIN chanx_right_in[0]
    PORT
      LAYER met3 ;
        RECT 96.000 54.440 100.000 55.040 ;
    END
  END chanx_right_in[0]
  PIN chanx_right_in[10]
    PORT
      LAYER met2 ;
        RECT 19.410 0.000 19.690 4.000 ;
    END
  END chanx_right_in[10]
  PIN chanx_right_in[1]
    PORT
      LAYER met3 ;
        RECT 96.000 37.440 100.000 38.040 ;
    END
  END chanx_right_in[1]
  PIN chanx_right_in[2]
    PORT
      LAYER met2 ;
        RECT 77.370 96.000 77.650 100.000 ;
    END
  END chanx_right_in[2]
  PIN chanx_right_in[3]
    PORT
      LAYER met2 ;
        RECT 77.370 0.000 77.650 4.000 ;
    END
  END chanx_right_in[3]
  PIN chanx_right_in[4]
    PORT
      LAYER met3 ;
        RECT 0.000 30.640 4.000 31.240 ;
    END
  END chanx_right_in[4]
  PIN chanx_right_in[5]
    PORT
      LAYER met3 ;
        RECT 0.000 44.240 4.000 44.840 ;
    END
  END chanx_right_in[5]
  PIN chanx_right_in[6]
    PORT
      LAYER met3 ;
        RECT 0.000 98.640 4.000 99.240 ;
    END
  END chanx_right_in[6]
  PIN chanx_right_in[7]
    PORT
      LAYER met3 ;
        RECT 96.000 17.040 100.000 17.640 ;
    END
  END chanx_right_in[7]
  PIN chanx_right_in[8]
    PORT
      LAYER met2 ;
        RECT 61.270 96.000 61.550 100.000 ;
    END
  END chanx_right_in[8]
  PIN chanx_right_in[9]
    PORT
      LAYER met3 ;
        RECT 0.000 61.240 4.000 61.840 ;
    END
  END chanx_right_in[9]
  PIN chanx_right_out[0]
    PORT
      LAYER met2 ;
        RECT 58.050 0.000 58.330 4.000 ;
    END
  END chanx_right_out[0]
  PIN chanx_right_out[10]
    PORT
      LAYER met3 ;
        RECT 96.000 23.840 100.000 24.440 ;
    END
  END chanx_right_out[10]
  PIN chanx_right_out[1]
    PORT
      LAYER met3 ;
        RECT 96.000 68.040 100.000 68.640 ;
    END
  END chanx_right_out[1]
  PIN chanx_right_out[2]
    PORT
      LAYER met2 ;
        RECT 3.310 96.000 3.590 100.000 ;
    END
  END chanx_right_out[2]
  PIN chanx_right_out[3]
    PORT
      LAYER met3 ;
        RECT 0.000 68.040 4.000 68.640 ;
    END
  END chanx_right_out[3]
  PIN chanx_right_out[4]
    PORT
      LAYER met3 ;
        RECT 96.000 91.840 100.000 92.440 ;
    END
  END chanx_right_out[4]
  PIN chanx_right_out[5]
    PORT
      LAYER met2 ;
        RECT 70.930 0.000 71.210 4.000 ;
    END
  END chanx_right_out[5]
  PIN chanx_right_out[6]
    PORT
      LAYER met2 ;
        RECT 87.030 0.000 87.310 4.000 ;
    END
  END chanx_right_out[6]
  PIN chanx_right_out[7]
    PORT
      LAYER met3 ;
        RECT 0.000 81.640 4.000 82.240 ;
    END
  END chanx_right_out[7]
  PIN chanx_right_out[8]
    PORT
      LAYER met3 ;
        RECT 96.000 0.040 100.000 0.640 ;
    END
  END chanx_right_out[8]
  PIN chanx_right_out[9]
    PORT
      LAYER met2 ;
        RECT 38.730 96.000 39.010 100.000 ;
    END
  END chanx_right_out[9]
  PIN chany_top_in[0]
    PORT
      LAYER met2 ;
        RECT 83.810 96.000 84.090 100.000 ;
    END
  END chany_top_in[0]
  PIN chany_top_in[10]
    PORT
      LAYER met3 ;
        RECT 0.000 13.640 4.000 14.240 ;
    END
  END chany_top_in[10]
  PIN chany_top_in[1]
    PORT
      LAYER met2 ;
        RECT 54.830 96.000 55.110 100.000 ;
    END
  END chany_top_in[1]
  PIN chany_top_in[2]
    PORT
      LAYER met3 ;
        RECT 0.000 20.440 4.000 21.040 ;
    END
  END chany_top_in[2]
  PIN chany_top_in[3]
    PORT
      LAYER met3 ;
        RECT 96.000 98.640 100.000 99.240 ;
    END
  END chany_top_in[3]
  PIN chany_top_in[4]
    PORT
      LAYER met3 ;
        RECT 96.000 78.240 100.000 78.840 ;
    END
  END chany_top_in[4]
  PIN chany_top_in[5]
    PORT
      LAYER met2 ;
        RECT 9.750 96.000 10.030 100.000 ;
    END
  END chany_top_in[5]
  PIN chany_top_in[6]
    PORT
      LAYER met2 ;
        RECT 67.710 96.000 67.990 100.000 ;
    END
  END chany_top_in[6]
  PIN chany_top_in[7]
    PORT
      LAYER met2 ;
        RECT 6.530 0.000 6.810 4.000 ;
    END
  END chany_top_in[7]
  PIN chany_top_in[8]
    PORT
      LAYER met2 ;
        RECT 0.090 0.000 0.370 4.000 ;
    END
  END chany_top_in[8]
  PIN chany_top_in[9]
    PORT
      LAYER met2 ;
        RECT 25.850 96.000 26.130 100.000 ;
    END
  END chany_top_in[9]
  PIN chany_top_out[0]
    PORT
      LAYER met3 ;
        RECT 96.000 85.040 100.000 85.640 ;
    END
  END chany_top_out[0]
  PIN chany_top_out[10]
    PORT
      LAYER met2 ;
        RECT 35.510 0.000 35.790 4.000 ;
    END
  END chany_top_out[10]
  PIN chany_top_out[1]
    PORT
      LAYER met3 ;
        RECT 96.000 61.240 100.000 61.840 ;
    END
  END chany_top_out[1]
  PIN chany_top_out[2]
    PORT
      LAYER met2 ;
        RECT 93.470 0.000 93.750 4.000 ;
    END
  END chany_top_out[2]
  PIN chany_top_out[3]
    PORT
      LAYER met2 ;
        RECT 48.390 96.000 48.670 100.000 ;
    END
  END chany_top_out[3]
  PIN chany_top_out[4]
    PORT
      LAYER met3 ;
        RECT 96.000 30.640 100.000 31.240 ;
    END
  END chany_top_out[4]
  PIN chany_top_out[5]
    PORT
      LAYER met2 ;
        RECT 12.970 0.000 13.250 4.000 ;
    END
  END chany_top_out[5]
  PIN chany_top_out[6]
    PORT
      LAYER met2 ;
        RECT 29.070 0.000 29.350 4.000 ;
    END
  END chany_top_out[6]
  PIN chany_top_out[7]
    PORT
      LAYER met2 ;
        RECT 41.950 0.000 42.230 4.000 ;
    END
  END chany_top_out[7]
  PIN chany_top_out[8]
    PORT
      LAYER met3 ;
        RECT 0.000 6.840 4.000 7.440 ;
    END
  END chany_top_out[8]
  PIN chany_top_out[9]
    PORT
      LAYER met2 ;
        RECT 48.390 0.000 48.670 4.000 ;
    END
  END chany_top_out[9]
  PIN prog_clk
    PORT
      LAYER met3 ;
        RECT 0.000 51.040 4.000 51.640 ;
    END
  END prog_clk
  PIN right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_
    PORT
      LAYER met2 ;
        RECT 90.250 96.000 90.530 100.000 ;
    END
  END right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_
  PIN right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_
    PORT
      LAYER met2 ;
        RECT 19.410 96.000 19.690 100.000 ;
    END
  END right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_
  PIN right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_
    PORT
      LAYER met2 ;
        RECT 32.290 96.000 32.570 100.000 ;
    END
  END right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_
  PIN right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_
    PORT
      LAYER met2 ;
        RECT 64.490 0.000 64.770 4.000 ;
    END
  END right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_
  PIN right_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_
    PORT
      LAYER met3 ;
        RECT 0.000 37.440 4.000 38.040 ;
    END
  END right_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_
  PIN right_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_
    PORT
      LAYER met3 ;
        RECT 0.000 91.840 4.000 92.440 ;
    END
  END right_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_
  PIN top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_
    PORT
      LAYER met3 ;
        RECT 96.000 47.640 100.000 48.240 ;
    END
  END top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_
  PIN vccd1
    PORT
      LAYER met4 ;
        RECT 82.400 10.640 84.000 87.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 60.205 10.640 61.805 87.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 38.010 10.640 39.610 87.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 15.815 10.640 17.415 87.280 ;
    END
  END vccd1
  PIN vssd1
    PORT
      LAYER met4 ;
        RECT 93.495 10.640 95.095 87.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 71.300 10.640 72.900 87.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 49.105 10.640 50.705 87.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 26.910 10.640 28.510 87.280 ;
    END
  END vssd1
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 94.300 87.125 ;
      LAYER met1 ;
        RECT 0.070 9.560 96.070 87.280 ;
      LAYER met2 ;
        RECT 0.100 95.720 3.030 99.125 ;
        RECT 3.870 95.720 9.470 99.125 ;
        RECT 10.310 95.720 19.130 99.125 ;
        RECT 19.970 95.720 25.570 99.125 ;
        RECT 26.410 95.720 32.010 99.125 ;
        RECT 32.850 95.720 38.450 99.125 ;
        RECT 39.290 95.720 48.110 99.125 ;
        RECT 48.950 95.720 54.550 99.125 ;
        RECT 55.390 95.720 60.990 99.125 ;
        RECT 61.830 95.720 67.430 99.125 ;
        RECT 68.270 95.720 77.090 99.125 ;
        RECT 77.930 95.720 83.530 99.125 ;
        RECT 84.370 95.720 89.970 99.125 ;
        RECT 90.810 95.720 96.050 99.125 ;
        RECT 0.100 4.280 96.050 95.720 ;
        RECT 0.650 0.155 6.250 4.280 ;
        RECT 7.090 0.155 12.690 4.280 ;
        RECT 13.530 0.155 19.130 4.280 ;
        RECT 19.970 0.155 28.790 4.280 ;
        RECT 29.630 0.155 35.230 4.280 ;
        RECT 36.070 0.155 41.670 4.280 ;
        RECT 42.510 0.155 48.110 4.280 ;
        RECT 48.950 0.155 57.770 4.280 ;
        RECT 58.610 0.155 64.210 4.280 ;
        RECT 65.050 0.155 70.650 4.280 ;
        RECT 71.490 0.155 77.090 4.280 ;
        RECT 77.930 0.155 86.750 4.280 ;
        RECT 87.590 0.155 93.190 4.280 ;
        RECT 94.030 0.155 96.050 4.280 ;
      LAYER met3 ;
        RECT 4.400 98.240 95.600 99.105 ;
        RECT 4.000 92.840 96.060 98.240 ;
        RECT 4.400 91.440 95.600 92.840 ;
        RECT 4.000 86.040 96.060 91.440 ;
        RECT 4.000 84.640 95.600 86.040 ;
        RECT 4.000 82.640 96.060 84.640 ;
        RECT 4.400 81.240 96.060 82.640 ;
        RECT 4.000 79.240 96.060 81.240 ;
        RECT 4.000 77.840 95.600 79.240 ;
        RECT 4.000 75.840 96.060 77.840 ;
        RECT 4.400 74.440 96.060 75.840 ;
        RECT 4.000 69.040 96.060 74.440 ;
        RECT 4.400 67.640 95.600 69.040 ;
        RECT 4.000 62.240 96.060 67.640 ;
        RECT 4.400 60.840 95.600 62.240 ;
        RECT 4.000 55.440 96.060 60.840 ;
        RECT 4.000 54.040 95.600 55.440 ;
        RECT 4.000 52.040 96.060 54.040 ;
        RECT 4.400 50.640 96.060 52.040 ;
        RECT 4.000 48.640 96.060 50.640 ;
        RECT 4.000 47.240 95.600 48.640 ;
        RECT 4.000 45.240 96.060 47.240 ;
        RECT 4.400 43.840 96.060 45.240 ;
        RECT 4.000 38.440 96.060 43.840 ;
        RECT 4.400 37.040 95.600 38.440 ;
        RECT 4.000 31.640 96.060 37.040 ;
        RECT 4.400 30.240 95.600 31.640 ;
        RECT 4.000 24.840 96.060 30.240 ;
        RECT 4.000 23.440 95.600 24.840 ;
        RECT 4.000 21.440 96.060 23.440 ;
        RECT 4.400 20.040 96.060 21.440 ;
        RECT 4.000 18.040 96.060 20.040 ;
        RECT 4.000 16.640 95.600 18.040 ;
        RECT 4.000 14.640 96.060 16.640 ;
        RECT 4.400 13.240 96.060 14.640 ;
        RECT 4.000 7.840 96.060 13.240 ;
        RECT 4.400 6.440 95.600 7.840 ;
        RECT 4.000 1.040 96.060 6.440 ;
        RECT 4.000 0.175 95.600 1.040 ;
  END
END sb_0__0_
END LIBRARY

