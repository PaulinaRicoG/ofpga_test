VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO cbx_1__0_
  CLASS BLOCK ;
  FOREIGN cbx_1__0_ ;
  ORIGIN 0.000 0.000 ;
  SIZE 100.000 BY 100.000 ;
  PIN bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_
    PORT
      LAYER met2 ;
        RECT 19.410 0.000 19.690 4.000 ;
    END
  END bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_
  PIN bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_
    PORT
      LAYER met3 ;
        RECT 0.000 61.240 4.000 61.840 ;
    END
  END bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_
  PIN bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_
    PORT
      LAYER met2 ;
        RECT 80.590 0.000 80.870 4.000 ;
    END
  END bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_
  PIN bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_
    PORT
      LAYER met2 ;
        RECT 6.530 96.000 6.810 100.000 ;
    END
  END bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_
  PIN bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_
    PORT
      LAYER met3 ;
        RECT 96.000 51.040 100.000 51.640 ;
    END
  END bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_
  PIN bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_
    PORT
      LAYER met2 ;
        RECT 74.150 0.000 74.430 4.000 ;
    END
  END bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_
  PIN ccff_head
    PORT
      LAYER met2 ;
        RECT 58.050 0.000 58.330 4.000 ;
    END
  END ccff_head
  PIN ccff_tail
    PORT
      LAYER met3 ;
        RECT 0.000 78.240 4.000 78.840 ;
    END
  END ccff_tail
  PIN chanx_left_in[0]
    PORT
      LAYER met3 ;
        RECT 0.000 98.640 4.000 99.240 ;
    END
  END chanx_left_in[0]
  PIN chanx_left_in[10]
    PORT
      LAYER met3 ;
        RECT 96.000 10.240 100.000 10.840 ;
    END
  END chanx_left_in[10]
  PIN chanx_left_in[1]
    PORT
      LAYER met2 ;
        RECT 64.490 96.000 64.770 100.000 ;
    END
  END chanx_left_in[1]
  PIN chanx_left_in[2]
    PORT
      LAYER met3 ;
        RECT 96.000 3.440 100.000 4.040 ;
    END
  END chanx_left_in[2]
  PIN chanx_left_in[3]
    PORT
      LAYER met2 ;
        RECT 80.590 96.000 80.870 100.000 ;
    END
  END chanx_left_in[3]
  PIN chanx_left_in[4]
    PORT
      LAYER met3 ;
        RECT 96.000 17.040 100.000 17.640 ;
    END
  END chanx_left_in[4]
  PIN chanx_left_in[5]
    PORT
      LAYER met2 ;
        RECT 12.970 96.000 13.250 100.000 ;
    END
  END chanx_left_in[5]
  PIN chanx_left_in[6]
    PORT
      LAYER met3 ;
        RECT 96.000 27.240 100.000 27.840 ;
    END
  END chanx_left_in[6]
  PIN chanx_left_in[7]
    PORT
      LAYER met3 ;
        RECT 0.000 68.040 4.000 68.640 ;
    END
  END chanx_left_in[7]
  PIN chanx_left_in[8]
    PORT
      LAYER met3 ;
        RECT 96.000 88.440 100.000 89.040 ;
    END
  END chanx_left_in[8]
  PIN chanx_left_in[9]
    PORT
      LAYER met3 ;
        RECT 0.000 30.640 4.000 31.240 ;
    END
  END chanx_left_in[9]
  PIN chanx_left_out[0]
    PORT
      LAYER met3 ;
        RECT 0.000 44.240 4.000 44.840 ;
    END
  END chanx_left_out[0]
  PIN chanx_left_out[10]
    PORT
      LAYER met3 ;
        RECT 0.000 85.040 4.000 85.640 ;
    END
  END chanx_left_out[10]
  PIN chanx_left_out[1]
    PORT
      LAYER met2 ;
        RECT 93.470 0.000 93.750 4.000 ;
    END
  END chanx_left_out[1]
  PIN chanx_left_out[2]
    PORT
      LAYER met3 ;
        RECT 0.000 54.440 4.000 55.040 ;
    END
  END chanx_left_out[2]
  PIN chanx_left_out[3]
    PORT
      LAYER met3 ;
        RECT 96.000 71.440 100.000 72.040 ;
    END
  END chanx_left_out[3]
  PIN chanx_left_out[4]
    PORT
      LAYER met3 ;
        RECT 0.000 13.640 4.000 14.240 ;
    END
  END chanx_left_out[4]
  PIN chanx_left_out[5]
    PORT
      LAYER met2 ;
        RECT 58.050 96.000 58.330 100.000 ;
    END
  END chanx_left_out[5]
  PIN chanx_left_out[6]
    PORT
      LAYER met3 ;
        RECT 0.000 20.440 4.000 21.040 ;
    END
  END chanx_left_out[6]
  PIN chanx_left_out[7]
    PORT
      LAYER met3 ;
        RECT 96.000 95.240 100.000 95.840 ;
    END
  END chanx_left_out[7]
  PIN chanx_left_out[8]
    PORT
      LAYER met2 ;
        RECT 41.950 96.000 42.230 100.000 ;
    END
  END chanx_left_out[8]
  PIN chanx_left_out[9]
    PORT
      LAYER met3 ;
        RECT 96.000 57.840 100.000 58.440 ;
    END
  END chanx_left_out[9]
  PIN chanx_right_in[0]
    PORT
      LAYER met2 ;
        RECT 70.930 96.000 71.210 100.000 ;
    END
  END chanx_right_in[0]
  PIN chanx_right_in[10]
    PORT
      LAYER met2 ;
        RECT 6.530 0.000 6.810 4.000 ;
    END
  END chanx_right_in[10]
  PIN chanx_right_in[1]
    PORT
      LAYER met2 ;
        RECT 0.090 0.000 0.370 4.000 ;
    END
  END chanx_right_in[1]
  PIN chanx_right_in[2]
    PORT
      LAYER met2 ;
        RECT 29.070 96.000 29.350 100.000 ;
    END
  END chanx_right_in[2]
  PIN chanx_right_in[3]
    PORT
      LAYER met3 ;
        RECT 96.000 81.640 100.000 82.240 ;
    END
  END chanx_right_in[3]
  PIN chanx_right_in[4]
    PORT
      LAYER met2 ;
        RECT 35.510 0.000 35.790 4.000 ;
    END
  END chanx_right_in[4]
  PIN chanx_right_in[5]
    PORT
      LAYER met3 ;
        RECT 96.000 64.640 100.000 65.240 ;
    END
  END chanx_right_in[5]
  PIN chanx_right_in[6]
    PORT
      LAYER met2 ;
        RECT 87.030 0.000 87.310 4.000 ;
    END
  END chanx_right_in[6]
  PIN chanx_right_in[7]
    PORT
      LAYER met2 ;
        RECT 51.610 96.000 51.890 100.000 ;
    END
  END chanx_right_in[7]
  PIN chanx_right_in[8]
    PORT
      LAYER met3 ;
        RECT 96.000 34.040 100.000 34.640 ;
    END
  END chanx_right_in[8]
  PIN chanx_right_in[9]
    PORT
      LAYER met2 ;
        RECT 12.970 0.000 13.250 4.000 ;
    END
  END chanx_right_in[9]
  PIN chanx_right_out[0]
    PORT
      LAYER met2 ;
        RECT 29.070 0.000 29.350 4.000 ;
    END
  END chanx_right_out[0]
  PIN chanx_right_out[10]
    PORT
      LAYER met2 ;
        RECT 41.950 0.000 42.230 4.000 ;
    END
  END chanx_right_out[10]
  PIN chanx_right_out[1]
    PORT
      LAYER met3 ;
        RECT 0.000 6.840 4.000 7.440 ;
    END
  END chanx_right_out[1]
  PIN chanx_right_out[2]
    PORT
      LAYER met2 ;
        RECT 51.610 0.000 51.890 4.000 ;
    END
  END chanx_right_out[2]
  PIN chanx_right_out[3]
    PORT
      LAYER met2 ;
        RECT 93.470 96.000 93.750 100.000 ;
    END
  END chanx_right_out[3]
  PIN chanx_right_out[4]
    PORT
      LAYER met2 ;
        RECT 87.030 96.000 87.310 100.000 ;
    END
  END chanx_right_out[4]
  PIN chanx_right_out[5]
    PORT
      LAYER met2 ;
        RECT 19.410 96.000 19.690 100.000 ;
    END
  END chanx_right_out[5]
  PIN chanx_right_out[6]
    PORT
      LAYER met2 ;
        RECT 35.510 96.000 35.790 100.000 ;
    END
  END chanx_right_out[6]
  PIN chanx_right_out[7]
    PORT
      LAYER met2 ;
        RECT 64.490 0.000 64.770 4.000 ;
    END
  END chanx_right_out[7]
  PIN chanx_right_out[8]
    PORT
      LAYER met3 ;
        RECT 0.000 37.440 4.000 38.040 ;
    END
  END chanx_right_out[8]
  PIN chanx_right_out[9]
    PORT
      LAYER met3 ;
        RECT 0.000 91.840 4.000 92.440 ;
    END
  END chanx_right_out[9]
  PIN prog_clk
    PORT
      LAYER met3 ;
        RECT 96.000 40.840 100.000 41.440 ;
    END
  END prog_clk
  PIN vccd1
    PORT
      LAYER met4 ;
        RECT 82.400 10.640 84.000 87.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 60.205 10.640 61.805 87.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 38.010 10.640 39.610 87.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 15.815 10.640 17.415 87.280 ;
    END
  END vccd1
  PIN vssd1
    PORT
      LAYER met4 ;
        RECT 93.495 10.640 95.095 87.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 71.300 10.640 72.900 87.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 49.105 10.640 50.705 87.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 26.910 10.640 28.510 87.280 ;
    END
  END vssd1
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 94.300 87.125 ;
      LAYER met1 ;
        RECT 0.070 10.240 96.070 87.280 ;
      LAYER met2 ;
        RECT 0.100 95.720 6.250 99.125 ;
        RECT 7.090 95.720 12.690 99.125 ;
        RECT 13.530 95.720 19.130 99.125 ;
        RECT 19.970 95.720 28.790 99.125 ;
        RECT 29.630 95.720 35.230 99.125 ;
        RECT 36.070 95.720 41.670 99.125 ;
        RECT 42.510 95.720 51.330 99.125 ;
        RECT 52.170 95.720 57.770 99.125 ;
        RECT 58.610 95.720 64.210 99.125 ;
        RECT 65.050 95.720 70.650 99.125 ;
        RECT 71.490 95.720 80.310 99.125 ;
        RECT 81.150 95.720 86.750 99.125 ;
        RECT 87.590 95.720 93.190 99.125 ;
        RECT 94.030 95.720 96.050 99.125 ;
        RECT 0.100 4.280 96.050 95.720 ;
        RECT 0.650 3.555 6.250 4.280 ;
        RECT 7.090 3.555 12.690 4.280 ;
        RECT 13.530 3.555 19.130 4.280 ;
        RECT 19.970 3.555 28.790 4.280 ;
        RECT 29.630 3.555 35.230 4.280 ;
        RECT 36.070 3.555 41.670 4.280 ;
        RECT 42.510 3.555 51.330 4.280 ;
        RECT 52.170 3.555 57.770 4.280 ;
        RECT 58.610 3.555 64.210 4.280 ;
        RECT 65.050 3.555 73.870 4.280 ;
        RECT 74.710 3.555 80.310 4.280 ;
        RECT 81.150 3.555 86.750 4.280 ;
        RECT 87.590 3.555 93.190 4.280 ;
        RECT 94.030 3.555 96.050 4.280 ;
      LAYER met3 ;
        RECT 4.400 98.240 96.075 99.105 ;
        RECT 4.000 96.240 96.075 98.240 ;
        RECT 4.000 94.840 95.600 96.240 ;
        RECT 4.000 92.840 96.075 94.840 ;
        RECT 4.400 91.440 96.075 92.840 ;
        RECT 4.000 89.440 96.075 91.440 ;
        RECT 4.000 88.040 95.600 89.440 ;
        RECT 4.000 86.040 96.075 88.040 ;
        RECT 4.400 84.640 96.075 86.040 ;
        RECT 4.000 82.640 96.075 84.640 ;
        RECT 4.000 81.240 95.600 82.640 ;
        RECT 4.000 79.240 96.075 81.240 ;
        RECT 4.400 77.840 96.075 79.240 ;
        RECT 4.000 72.440 96.075 77.840 ;
        RECT 4.000 71.040 95.600 72.440 ;
        RECT 4.000 69.040 96.075 71.040 ;
        RECT 4.400 67.640 96.075 69.040 ;
        RECT 4.000 65.640 96.075 67.640 ;
        RECT 4.000 64.240 95.600 65.640 ;
        RECT 4.000 62.240 96.075 64.240 ;
        RECT 4.400 60.840 96.075 62.240 ;
        RECT 4.000 58.840 96.075 60.840 ;
        RECT 4.000 57.440 95.600 58.840 ;
        RECT 4.000 55.440 96.075 57.440 ;
        RECT 4.400 54.040 96.075 55.440 ;
        RECT 4.000 52.040 96.075 54.040 ;
        RECT 4.000 50.640 95.600 52.040 ;
        RECT 4.000 45.240 96.075 50.640 ;
        RECT 4.400 43.840 96.075 45.240 ;
        RECT 4.000 41.840 96.075 43.840 ;
        RECT 4.000 40.440 95.600 41.840 ;
        RECT 4.000 38.440 96.075 40.440 ;
        RECT 4.400 37.040 96.075 38.440 ;
        RECT 4.000 35.040 96.075 37.040 ;
        RECT 4.000 33.640 95.600 35.040 ;
        RECT 4.000 31.640 96.075 33.640 ;
        RECT 4.400 30.240 96.075 31.640 ;
        RECT 4.000 28.240 96.075 30.240 ;
        RECT 4.000 26.840 95.600 28.240 ;
        RECT 4.000 21.440 96.075 26.840 ;
        RECT 4.400 20.040 96.075 21.440 ;
        RECT 4.000 18.040 96.075 20.040 ;
        RECT 4.000 16.640 95.600 18.040 ;
        RECT 4.000 14.640 96.075 16.640 ;
        RECT 4.400 13.240 96.075 14.640 ;
        RECT 4.000 11.240 96.075 13.240 ;
        RECT 4.000 9.840 95.600 11.240 ;
        RECT 4.000 7.840 96.075 9.840 ;
        RECT 4.400 6.440 96.075 7.840 ;
        RECT 4.000 4.440 96.075 6.440 ;
        RECT 4.000 3.575 95.600 4.440 ;
      LAYER met4 ;
        RECT 84.935 27.375 85.265 36.545 ;
  END
END cbx_1__0_
END LIBRARY

