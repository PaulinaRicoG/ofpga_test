VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sb_1__4_
  CLASS BLOCK ;
  FOREIGN sb_1__4_ ;
  ORIGIN 0.000 0.000 ;
  SIZE 100.000 BY 100.000 ;
  PIN bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_
    PORT
      LAYER met2 ;
        RECT 32.290 96.000 32.570 100.000 ;
    END
  END bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_
  PIN bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_
    PORT
      LAYER met2 ;
        RECT 64.490 96.000 64.770 100.000 ;
    END
  END bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_
  PIN bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_12_
    PORT
      LAYER met2 ;
        RECT 9.750 0.000 10.030 4.000 ;
    END
  END bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_12_
  PIN bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_13_
    PORT
      LAYER met3 ;
        RECT 0.000 10.240 4.000 10.840 ;
    END
  END bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_13_
  PIN bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_14_
    PORT
      LAYER met3 ;
        RECT 96.000 0.040 100.000 0.640 ;
    END
  END bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_14_
  PIN bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_
    PORT
      LAYER met3 ;
        RECT 96.000 34.040 100.000 34.640 ;
    END
  END bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_
  PIN bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_
    PORT
      LAYER met2 ;
        RECT 87.030 96.000 87.310 100.000 ;
    END
  END bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_
  PIN ccff_head
    PORT
      LAYER met3 ;
        RECT 96.000 51.040 100.000 51.640 ;
    END
  END ccff_head
  PIN ccff_tail
    PORT
      LAYER met3 ;
        RECT 96.000 81.640 100.000 82.240 ;
    END
  END ccff_tail
  PIN chanx_left_in[0]
    PORT
      LAYER met3 ;
        RECT 0.000 81.640 4.000 82.240 ;
    END
  END chanx_left_in[0]
  PIN chanx_left_in[10]
    PORT
      LAYER met2 ;
        RECT 35.510 0.000 35.790 4.000 ;
    END
  END chanx_left_in[10]
  PIN chanx_left_in[1]
    PORT
      LAYER met2 ;
        RECT 48.390 96.000 48.670 100.000 ;
    END
  END chanx_left_in[1]
  PIN chanx_left_in[2]
    PORT
      LAYER met3 ;
        RECT 96.000 68.040 100.000 68.640 ;
    END
  END chanx_left_in[2]
  PIN chanx_left_in[3]
    PORT
      LAYER met2 ;
        RECT 93.470 0.000 93.750 4.000 ;
    END
  END chanx_left_in[3]
  PIN chanx_left_in[4]
    PORT
      LAYER met3 ;
        RECT 0.000 74.840 4.000 75.440 ;
    END
  END chanx_left_in[4]
  PIN chanx_left_in[5]
    PORT
      LAYER met2 ;
        RECT 3.310 96.000 3.590 100.000 ;
    END
  END chanx_left_in[5]
  PIN chanx_left_in[6]
    PORT
      LAYER met2 ;
        RECT 38.730 96.000 39.010 100.000 ;
    END
  END chanx_left_in[6]
  PIN chanx_left_in[7]
    PORT
      LAYER met3 ;
        RECT 0.000 20.440 4.000 21.040 ;
    END
  END chanx_left_in[7]
  PIN chanx_left_in[8]
    PORT
      LAYER met3 ;
        RECT 96.000 88.440 100.000 89.040 ;
    END
  END chanx_left_in[8]
  PIN chanx_left_in[9]
    PORT
      LAYER met3 ;
        RECT 96.000 20.440 100.000 21.040 ;
    END
  END chanx_left_in[9]
  PIN chanx_left_out[0]
    PORT
      LAYER met2 ;
        RECT 67.710 96.000 67.990 100.000 ;
    END
  END chanx_left_out[0]
  PIN chanx_left_out[10]
    PORT
      LAYER met2 ;
        RECT 22.630 0.000 22.910 4.000 ;
    END
  END chanx_left_out[10]
  PIN chanx_left_out[1]
    PORT
      LAYER met3 ;
        RECT 96.000 74.840 100.000 75.440 ;
    END
  END chanx_left_out[1]
  PIN chanx_left_out[2]
    PORT
      LAYER met2 ;
        RECT 77.370 0.000 77.650 4.000 ;
    END
  END chanx_left_out[2]
  PIN chanx_left_out[3]
    PORT
      LAYER met2 ;
        RECT 90.250 96.000 90.530 100.000 ;
    END
  END chanx_left_out[3]
  PIN chanx_left_out[4]
    PORT
      LAYER met3 ;
        RECT 96.000 13.640 100.000 14.240 ;
    END
  END chanx_left_out[4]
  PIN chanx_left_out[5]
    PORT
      LAYER met2 ;
        RECT 58.050 96.000 58.330 100.000 ;
    END
  END chanx_left_out[5]
  PIN chanx_left_out[6]
    PORT
      LAYER met3 ;
        RECT 96.000 78.240 100.000 78.840 ;
    END
  END chanx_left_out[6]
  PIN chanx_left_out[7]
    PORT
      LAYER met3 ;
        RECT 0.000 98.640 4.000 99.240 ;
    END
  END chanx_left_out[7]
  PIN chanx_left_out[8]
    PORT
      LAYER met3 ;
        RECT 0.000 3.440 4.000 4.040 ;
    END
  END chanx_left_out[8]
  PIN chanx_left_out[9]
    PORT
      LAYER met3 ;
        RECT 0.000 47.640 4.000 48.240 ;
    END
  END chanx_left_out[9]
  PIN chanx_right_in[0]
    PORT
      LAYER met2 ;
        RECT 19.410 0.000 19.690 4.000 ;
    END
  END chanx_right_in[0]
  PIN chanx_right_in[10]
    PORT
      LAYER met2 ;
        RECT 45.170 96.000 45.450 100.000 ;
    END
  END chanx_right_in[10]
  PIN chanx_right_in[1]
    PORT
      LAYER met3 ;
        RECT 96.000 64.640 100.000 65.240 ;
    END
  END chanx_right_in[1]
  PIN chanx_right_in[2]
    PORT
      LAYER met3 ;
        RECT 96.000 23.840 100.000 24.440 ;
    END
  END chanx_right_in[2]
  PIN chanx_right_in[3]
    PORT
      LAYER met2 ;
        RECT 61.270 96.000 61.550 100.000 ;
    END
  END chanx_right_in[3]
  PIN chanx_right_in[4]
    PORT
      LAYER met3 ;
        RECT 0.000 6.840 4.000 7.440 ;
    END
  END chanx_right_in[4]
  PIN chanx_right_in[5]
    PORT
      LAYER met2 ;
        RECT 90.250 0.000 90.530 4.000 ;
    END
  END chanx_right_in[5]
  PIN chanx_right_in[6]
    PORT
      LAYER met2 ;
        RECT 35.510 96.000 35.790 100.000 ;
    END
  END chanx_right_in[6]
  PIN chanx_right_in[7]
    PORT
      LAYER met3 ;
        RECT 96.000 91.840 100.000 92.440 ;
    END
  END chanx_right_in[7]
  PIN chanx_right_in[8]
    PORT
      LAYER met2 ;
        RECT 61.270 0.000 61.550 4.000 ;
    END
  END chanx_right_in[8]
  PIN chanx_right_in[9]
    PORT
      LAYER met3 ;
        RECT 0.000 51.040 4.000 51.640 ;
    END
  END chanx_right_in[9]
  PIN chanx_right_out[0]
    PORT
      LAYER met3 ;
        RECT 0.000 68.040 4.000 68.640 ;
    END
  END chanx_right_out[0]
  PIN chanx_right_out[10]
    PORT
      LAYER met3 ;
        RECT 96.000 44.240 100.000 44.840 ;
    END
  END chanx_right_out[10]
  PIN chanx_right_out[1]
    PORT
      LAYER met3 ;
        RECT 0.000 95.240 4.000 95.840 ;
    END
  END chanx_right_out[1]
  PIN chanx_right_out[2]
    PORT
      LAYER met2 ;
        RECT 80.590 0.000 80.870 4.000 ;
    END
  END chanx_right_out[2]
  PIN chanx_right_out[3]
    PORT
      LAYER met2 ;
        RECT 38.730 0.000 39.010 4.000 ;
    END
  END chanx_right_out[3]
  PIN chanx_right_out[4]
    PORT
      LAYER met2 ;
        RECT 70.930 0.000 71.210 4.000 ;
    END
  END chanx_right_out[4]
  PIN chanx_right_out[5]
    PORT
      LAYER met2 ;
        RECT 96.690 96.000 96.970 100.000 ;
    END
  END chanx_right_out[5]
  PIN chanx_right_out[6]
    PORT
      LAYER met2 ;
        RECT 16.190 96.000 16.470 100.000 ;
    END
  END chanx_right_out[6]
  PIN chanx_right_out[7]
    PORT
      LAYER met2 ;
        RECT 6.530 0.000 6.810 4.000 ;
    END
  END chanx_right_out[7]
  PIN chanx_right_out[8]
    PORT
      LAYER met2 ;
        RECT 29.070 0.000 29.350 4.000 ;
    END
  END chanx_right_out[8]
  PIN chanx_right_out[9]
    PORT
      LAYER met2 ;
        RECT 87.030 0.000 87.310 4.000 ;
    END
  END chanx_right_out[9]
  PIN chany_bottom_in[0]
    PORT
      LAYER met3 ;
        RECT 96.000 37.440 100.000 38.040 ;
    END
  END chany_bottom_in[0]
  PIN chany_bottom_in[10]
    PORT
      LAYER met3 ;
        RECT 96.000 17.040 100.000 17.640 ;
    END
  END chany_bottom_in[10]
  PIN chany_bottom_in[1]
    PORT
      LAYER met3 ;
        RECT 0.000 17.040 4.000 17.640 ;
    END
  END chany_bottom_in[1]
  PIN chany_bottom_in[2]
    PORT
      LAYER met3 ;
        RECT 0.000 91.840 4.000 92.440 ;
    END
  END chany_bottom_in[2]
  PIN chany_bottom_in[3]
    PORT
      LAYER met3 ;
        RECT 96.000 3.440 100.000 4.040 ;
    END
  END chany_bottom_in[3]
  PIN chany_bottom_in[4]
    PORT
      LAYER met2 ;
        RECT 19.410 96.000 19.690 100.000 ;
    END
  END chany_bottom_in[4]
  PIN chany_bottom_in[5]
    PORT
      LAYER met3 ;
        RECT 96.000 30.640 100.000 31.240 ;
    END
  END chany_bottom_in[5]
  PIN chany_bottom_in[6]
    PORT
      LAYER met3 ;
        RECT 0.000 61.240 4.000 61.840 ;
    END
  END chany_bottom_in[6]
  PIN chany_bottom_in[7]
    PORT
      LAYER met2 ;
        RECT 74.150 0.000 74.430 4.000 ;
    END
  END chany_bottom_in[7]
  PIN chany_bottom_in[8]
    PORT
      LAYER met3 ;
        RECT 96.000 61.240 100.000 61.840 ;
    END
  END chany_bottom_in[8]
  PIN chany_bottom_in[9]
    PORT
      LAYER met3 ;
        RECT 0.000 78.240 4.000 78.840 ;
    END
  END chany_bottom_in[9]
  PIN chany_bottom_out[0]
    PORT
      LAYER met2 ;
        RECT 9.750 96.000 10.030 100.000 ;
    END
  END chany_bottom_out[0]
  PIN chany_bottom_out[10]
    PORT
      LAYER met2 ;
        RECT 48.390 0.000 48.670 4.000 ;
    END
  END chany_bottom_out[10]
  PIN chany_bottom_out[1]
    PORT
      LAYER met2 ;
        RECT 0.090 0.000 0.370 4.000 ;
    END
  END chany_bottom_out[1]
  PIN chany_bottom_out[2]
    PORT
      LAYER met2 ;
        RECT 58.050 0.000 58.330 4.000 ;
    END
  END chany_bottom_out[2]
  PIN chany_bottom_out[3]
    PORT
      LAYER met2 ;
        RECT 25.850 96.000 26.130 100.000 ;
    END
  END chany_bottom_out[3]
  PIN chany_bottom_out[4]
    PORT
      LAYER met2 ;
        RECT 51.610 96.000 51.890 100.000 ;
    END
  END chany_bottom_out[4]
  PIN chany_bottom_out[5]
    PORT
      LAYER met3 ;
        RECT 0.000 34.040 4.000 34.640 ;
    END
  END chany_bottom_out[5]
  PIN chany_bottom_out[6]
    PORT
      LAYER met3 ;
        RECT 0.000 64.640 4.000 65.240 ;
    END
  END chany_bottom_out[6]
  PIN chany_bottom_out[7]
    PORT
      LAYER met3 ;
        RECT 0.000 54.440 4.000 55.040 ;
    END
  END chany_bottom_out[7]
  PIN chany_bottom_out[8]
    PORT
      LAYER met2 ;
        RECT 3.310 0.000 3.590 4.000 ;
    END
  END chany_bottom_out[8]
  PIN chany_bottom_out[9]
    PORT
      LAYER met2 ;
        RECT 93.470 96.000 93.750 100.000 ;
    END
  END chany_bottom_out[9]
  PIN left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_
    PORT
      LAYER met2 ;
        RECT 74.150 96.000 74.430 100.000 ;
    END
  END left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_
  PIN left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_
    PORT
      LAYER met2 ;
        RECT 45.170 0.000 45.450 4.000 ;
    END
  END left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_
  PIN left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_
    PORT
      LAYER met3 ;
        RECT 96.000 95.240 100.000 95.840 ;
    END
  END left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_
  PIN left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_
    PORT
      LAYER met3 ;
        RECT 96.000 6.840 100.000 7.440 ;
    END
  END left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_
  PIN left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_
    PORT
      LAYER met3 ;
        RECT 0.000 23.840 4.000 24.440 ;
    END
  END left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_
  PIN left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_
    PORT
      LAYER met3 ;
        RECT 0.000 40.840 4.000 41.440 ;
    END
  END left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_
  PIN left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_
    PORT
      LAYER met2 ;
        RECT 16.190 0.000 16.470 4.000 ;
    END
  END left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_
  PIN left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_
    PORT
      LAYER met2 ;
        RECT 32.290 0.000 32.570 4.000 ;
    END
  END left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_
  PIN left_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_
    PORT
      LAYER met3 ;
        RECT 0.000 37.440 4.000 38.040 ;
    END
  END left_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_
  PIN prog_clk
    PORT
      LAYER met3 ;
        RECT 96.000 57.840 100.000 58.440 ;
    END
  END prog_clk
  PIN right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_
    PORT
      LAYER met2 ;
        RECT 51.610 0.000 51.890 4.000 ;
    END
  END right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_
  PIN right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_
    PORT
      LAYER met2 ;
        RECT 80.590 96.000 80.870 100.000 ;
    END
  END right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_
  PIN right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_
    PORT
      LAYER met2 ;
        RECT 77.370 96.000 77.650 100.000 ;
    END
  END right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_
  PIN right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_
    PORT
      LAYER met2 ;
        RECT 6.530 96.000 6.810 100.000 ;
    END
  END right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_
  PIN right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_
    PORT
      LAYER met2 ;
        RECT 22.630 96.000 22.910 100.000 ;
    END
  END right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_
  PIN right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_
    PORT
      LAYER met2 ;
        RECT 64.490 0.000 64.770 4.000 ;
    END
  END right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_
  PIN right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_
    PORT
      LAYER met3 ;
        RECT 0.000 30.640 4.000 31.240 ;
    END
  END right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_
  PIN right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_
    PORT
      LAYER met3 ;
        RECT 0.000 85.040 4.000 85.640 ;
    END
  END right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_
  PIN right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_
    PORT
      LAYER met3 ;
        RECT 96.000 47.640 100.000 48.240 ;
    END
  END right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_
  PIN vccd1
    PORT
      LAYER met4 ;
        RECT 82.400 10.640 84.000 87.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 60.205 10.640 61.805 87.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 38.010 10.640 39.610 87.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 15.815 10.640 17.415 87.280 ;
    END
  END vccd1
  PIN vssd1
    PORT
      LAYER met4 ;
        RECT 93.495 10.640 95.095 87.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 71.300 10.640 72.900 87.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 49.105 10.640 50.705 87.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 26.910 10.640 28.510 87.280 ;
    END
  END vssd1
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 94.300 87.125 ;
      LAYER met1 ;
        RECT 0.070 10.240 96.990 88.020 ;
      LAYER met2 ;
        RECT 0.100 95.720 3.030 99.125 ;
        RECT 3.870 95.720 6.250 99.125 ;
        RECT 7.090 95.720 9.470 99.125 ;
        RECT 10.310 95.720 15.910 99.125 ;
        RECT 16.750 95.720 19.130 99.125 ;
        RECT 19.970 95.720 22.350 99.125 ;
        RECT 23.190 95.720 25.570 99.125 ;
        RECT 26.410 95.720 32.010 99.125 ;
        RECT 32.850 95.720 35.230 99.125 ;
        RECT 36.070 95.720 38.450 99.125 ;
        RECT 39.290 95.720 44.890 99.125 ;
        RECT 45.730 95.720 48.110 99.125 ;
        RECT 48.950 95.720 51.330 99.125 ;
        RECT 52.170 95.720 57.770 99.125 ;
        RECT 58.610 95.720 60.990 99.125 ;
        RECT 61.830 95.720 64.210 99.125 ;
        RECT 65.050 95.720 67.430 99.125 ;
        RECT 68.270 95.720 73.870 99.125 ;
        RECT 74.710 95.720 77.090 99.125 ;
        RECT 77.930 95.720 80.310 99.125 ;
        RECT 81.150 95.720 86.750 99.125 ;
        RECT 87.590 95.720 89.970 99.125 ;
        RECT 90.810 95.720 93.190 99.125 ;
        RECT 94.030 95.720 96.410 99.125 ;
        RECT 0.100 4.280 96.960 95.720 ;
        RECT 0.650 0.155 3.030 4.280 ;
        RECT 3.870 0.155 6.250 4.280 ;
        RECT 7.090 0.155 9.470 4.280 ;
        RECT 10.310 0.155 15.910 4.280 ;
        RECT 16.750 0.155 19.130 4.280 ;
        RECT 19.970 0.155 22.350 4.280 ;
        RECT 23.190 0.155 28.790 4.280 ;
        RECT 29.630 0.155 32.010 4.280 ;
        RECT 32.850 0.155 35.230 4.280 ;
        RECT 36.070 0.155 38.450 4.280 ;
        RECT 39.290 0.155 44.890 4.280 ;
        RECT 45.730 0.155 48.110 4.280 ;
        RECT 48.950 0.155 51.330 4.280 ;
        RECT 52.170 0.155 57.770 4.280 ;
        RECT 58.610 0.155 60.990 4.280 ;
        RECT 61.830 0.155 64.210 4.280 ;
        RECT 65.050 0.155 70.650 4.280 ;
        RECT 71.490 0.155 73.870 4.280 ;
        RECT 74.710 0.155 77.090 4.280 ;
        RECT 77.930 0.155 80.310 4.280 ;
        RECT 81.150 0.155 86.750 4.280 ;
        RECT 87.590 0.155 89.970 4.280 ;
        RECT 90.810 0.155 93.190 4.280 ;
        RECT 94.030 0.155 96.960 4.280 ;
      LAYER met3 ;
        RECT 4.400 98.240 97.210 99.105 ;
        RECT 4.000 96.240 97.210 98.240 ;
        RECT 4.400 94.840 95.600 96.240 ;
        RECT 4.000 92.840 97.210 94.840 ;
        RECT 4.400 91.440 95.600 92.840 ;
        RECT 4.000 89.440 97.210 91.440 ;
        RECT 4.000 88.040 95.600 89.440 ;
        RECT 4.000 86.040 97.210 88.040 ;
        RECT 4.400 84.640 97.210 86.040 ;
        RECT 4.000 82.640 97.210 84.640 ;
        RECT 4.400 81.240 95.600 82.640 ;
        RECT 4.000 79.240 97.210 81.240 ;
        RECT 4.400 77.840 95.600 79.240 ;
        RECT 4.000 75.840 97.210 77.840 ;
        RECT 4.400 74.440 95.600 75.840 ;
        RECT 4.000 69.040 97.210 74.440 ;
        RECT 4.400 67.640 95.600 69.040 ;
        RECT 4.000 65.640 97.210 67.640 ;
        RECT 4.400 64.240 95.600 65.640 ;
        RECT 4.000 62.240 97.210 64.240 ;
        RECT 4.400 60.840 95.600 62.240 ;
        RECT 4.000 58.840 97.210 60.840 ;
        RECT 4.000 57.440 95.600 58.840 ;
        RECT 4.000 55.440 97.210 57.440 ;
        RECT 4.400 54.040 97.210 55.440 ;
        RECT 4.000 52.040 97.210 54.040 ;
        RECT 4.400 50.640 95.600 52.040 ;
        RECT 4.000 48.640 97.210 50.640 ;
        RECT 4.400 47.240 95.600 48.640 ;
        RECT 4.000 45.240 97.210 47.240 ;
        RECT 4.000 43.840 95.600 45.240 ;
        RECT 4.000 41.840 97.210 43.840 ;
        RECT 4.400 40.440 97.210 41.840 ;
        RECT 4.000 38.440 97.210 40.440 ;
        RECT 4.400 37.040 95.600 38.440 ;
        RECT 4.000 35.040 97.210 37.040 ;
        RECT 4.400 33.640 95.600 35.040 ;
        RECT 4.000 31.640 97.210 33.640 ;
        RECT 4.400 30.240 95.600 31.640 ;
        RECT 4.000 24.840 97.210 30.240 ;
        RECT 4.400 23.440 95.600 24.840 ;
        RECT 4.000 21.440 97.210 23.440 ;
        RECT 4.400 20.040 95.600 21.440 ;
        RECT 4.000 18.040 97.210 20.040 ;
        RECT 4.400 16.640 95.600 18.040 ;
        RECT 4.000 14.640 97.210 16.640 ;
        RECT 4.000 13.240 95.600 14.640 ;
        RECT 4.000 11.240 97.210 13.240 ;
        RECT 4.400 9.840 97.210 11.240 ;
        RECT 4.000 7.840 97.210 9.840 ;
        RECT 4.400 6.440 95.600 7.840 ;
        RECT 4.000 4.440 97.210 6.440 ;
        RECT 4.400 3.040 95.600 4.440 ;
        RECT 4.000 1.040 97.210 3.040 ;
        RECT 4.000 0.175 95.600 1.040 ;
      LAYER met4 ;
        RECT 62.855 13.095 70.900 80.065 ;
        RECT 73.300 13.095 82.000 80.065 ;
        RECT 84.400 13.095 90.785 80.065 ;
  END
END sb_1__4_
END LIBRARY

