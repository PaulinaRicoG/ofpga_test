VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sb_0__4_
  CLASS BLOCK ;
  FOREIGN sb_0__4_ ;
  ORIGIN 0.000 0.000 ;
  SIZE 100.000 BY 100.000 ;
  PIN bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_
    PORT
      LAYER met2 ;
        RECT 54.830 0.000 55.110 4.000 ;
    END
  END bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_
  PIN ccff_head
    PORT
      LAYER met3 ;
        RECT 96.000 17.040 100.000 17.640 ;
    END
  END ccff_head
  PIN ccff_tail
    PORT
      LAYER met3 ;
        RECT 96.000 3.440 100.000 4.040 ;
    END
  END ccff_tail
  PIN chanx_right_in[0]
    PORT
      LAYER met2 ;
        RECT 6.530 0.000 6.810 4.000 ;
    END
  END chanx_right_in[0]
  PIN chanx_right_in[10]
    PORT
      LAYER met2 ;
        RECT 61.270 96.000 61.550 100.000 ;
    END
  END chanx_right_in[10]
  PIN chanx_right_in[1]
    PORT
      LAYER met3 ;
        RECT 96.000 54.440 100.000 55.040 ;
    END
  END chanx_right_in[1]
  PIN chanx_right_in[2]
    PORT
      LAYER met3 ;
        RECT 96.000 23.840 100.000 24.440 ;
    END
  END chanx_right_in[2]
  PIN chanx_right_in[3]
    PORT
      LAYER met2 ;
        RECT 87.030 0.000 87.310 4.000 ;
    END
  END chanx_right_in[3]
  PIN chanx_right_in[4]
    PORT
      LAYER met3 ;
        RECT 96.000 74.840 100.000 75.440 ;
    END
  END chanx_right_in[4]
  PIN chanx_right_in[5]
    PORT
      LAYER met3 ;
        RECT 96.000 61.240 100.000 61.840 ;
    END
  END chanx_right_in[5]
  PIN chanx_right_in[6]
    PORT
      LAYER met3 ;
        RECT 96.000 81.640 100.000 82.240 ;
    END
  END chanx_right_in[6]
  PIN chanx_right_in[7]
    PORT
      LAYER met2 ;
        RECT 74.150 0.000 74.430 4.000 ;
    END
  END chanx_right_in[7]
  PIN chanx_right_in[8]
    PORT
      LAYER met2 ;
        RECT 19.410 0.000 19.690 4.000 ;
    END
  END chanx_right_in[8]
  PIN chanx_right_in[9]
    PORT
      LAYER met3 ;
        RECT 96.000 30.640 100.000 31.240 ;
    END
  END chanx_right_in[9]
  PIN chanx_right_out[0]
    PORT
      LAYER met2 ;
        RECT 54.830 96.000 55.110 100.000 ;
    END
  END chanx_right_out[0]
  PIN chanx_right_out[10]
    PORT
      LAYER met2 ;
        RECT 80.590 96.000 80.870 100.000 ;
    END
  END chanx_right_out[10]
  PIN chanx_right_out[1]
    PORT
      LAYER met2 ;
        RECT 67.710 0.000 67.990 4.000 ;
    END
  END chanx_right_out[1]
  PIN chanx_right_out[2]
    PORT
      LAYER met3 ;
        RECT 0.000 98.640 4.000 99.240 ;
    END
  END chanx_right_out[2]
  PIN chanx_right_out[3]
    PORT
      LAYER met3 ;
        RECT 96.000 95.240 100.000 95.840 ;
    END
  END chanx_right_out[3]
  PIN chanx_right_out[4]
    PORT
      LAYER met3 ;
        RECT 0.000 71.440 4.000 72.040 ;
    END
  END chanx_right_out[4]
  PIN chanx_right_out[5]
    PORT
      LAYER met3 ;
        RECT 0.000 27.240 4.000 27.840 ;
    END
  END chanx_right_out[5]
  PIN chanx_right_out[6]
    PORT
      LAYER met3 ;
        RECT 0.000 57.840 4.000 58.440 ;
    END
  END chanx_right_out[6]
  PIN chanx_right_out[7]
    PORT
      LAYER met2 ;
        RECT 80.590 0.000 80.870 4.000 ;
    END
  END chanx_right_out[7]
  PIN chanx_right_out[8]
    PORT
      LAYER met2 ;
        RECT 12.970 96.000 13.250 100.000 ;
    END
  END chanx_right_out[8]
  PIN chanx_right_out[9]
    PORT
      LAYER met3 ;
        RECT 0.000 78.240 4.000 78.840 ;
    END
  END chanx_right_out[9]
  PIN chany_bottom_in[0]
    PORT
      LAYER met3 ;
        RECT 96.000 10.240 100.000 10.840 ;
    END
  END chany_bottom_in[0]
  PIN chany_bottom_in[10]
    PORT
      LAYER met3 ;
        RECT 0.000 85.040 4.000 85.640 ;
    END
  END chany_bottom_in[10]
  PIN chany_bottom_in[1]
    PORT
      LAYER met2 ;
        RECT 74.150 96.000 74.430 100.000 ;
    END
  END chany_bottom_in[1]
  PIN chany_bottom_in[2]
    PORT
      LAYER met2 ;
        RECT 25.850 96.000 26.130 100.000 ;
    END
  END chany_bottom_in[2]
  PIN chany_bottom_in[3]
    PORT
      LAYER met2 ;
        RECT 45.170 96.000 45.450 100.000 ;
    END
  END chany_bottom_in[3]
  PIN chany_bottom_in[4]
    PORT
      LAYER met2 ;
        RECT 38.730 0.000 39.010 4.000 ;
    END
  END chany_bottom_in[4]
  PIN chany_bottom_in[5]
    PORT
      LAYER met3 ;
        RECT 0.000 47.640 4.000 48.240 ;
    END
  END chany_bottom_in[5]
  PIN chany_bottom_in[6]
    PORT
      LAYER met3 ;
        RECT 0.000 20.440 4.000 21.040 ;
    END
  END chany_bottom_in[6]
  PIN chany_bottom_in[7]
    PORT
      LAYER met2 ;
        RECT 6.530 96.000 6.810 100.000 ;
    END
  END chany_bottom_in[7]
  PIN chany_bottom_in[8]
    PORT
      LAYER met2 ;
        RECT 67.710 96.000 67.990 100.000 ;
    END
  END chany_bottom_in[8]
  PIN chany_bottom_in[9]
    PORT
      LAYER met3 ;
        RECT 0.000 13.640 4.000 14.240 ;
    END
  END chany_bottom_in[9]
  PIN chany_bottom_out[0]
    PORT
      LAYER met2 ;
        RECT 0.090 0.000 0.370 4.000 ;
    END
  END chany_bottom_out[0]
  PIN chany_bottom_out[10]
    PORT
      LAYER met3 ;
        RECT 0.000 40.840 4.000 41.440 ;
    END
  END chany_bottom_out[10]
  PIN chany_bottom_out[1]
    PORT
      LAYER met3 ;
        RECT 96.000 88.440 100.000 89.040 ;
    END
  END chany_bottom_out[1]
  PIN chany_bottom_out[2]
    PORT
      LAYER met2 ;
        RECT 32.290 0.000 32.570 4.000 ;
    END
  END chany_bottom_out[2]
  PIN chany_bottom_out[3]
    PORT
      LAYER met3 ;
        RECT 96.000 68.040 100.000 68.640 ;
    END
  END chany_bottom_out[3]
  PIN chany_bottom_out[4]
    PORT
      LAYER met2 ;
        RECT 93.470 0.000 93.750 4.000 ;
    END
  END chany_bottom_out[4]
  PIN chany_bottom_out[5]
    PORT
      LAYER met2 ;
        RECT 38.730 96.000 39.010 100.000 ;
    END
  END chany_bottom_out[5]
  PIN chany_bottom_out[6]
    PORT
      LAYER met3 ;
        RECT 96.000 37.440 100.000 38.040 ;
    END
  END chany_bottom_out[6]
  PIN chany_bottom_out[7]
    PORT
      LAYER met2 ;
        RECT 12.970 0.000 13.250 4.000 ;
    END
  END chany_bottom_out[7]
  PIN chany_bottom_out[8]
    PORT
      LAYER met2 ;
        RECT 25.850 0.000 26.130 4.000 ;
    END
  END chany_bottom_out[8]
  PIN chany_bottom_out[9]
    PORT
      LAYER met3 ;
        RECT 0.000 64.640 4.000 65.240 ;
    END
  END chany_bottom_out[9]
  PIN prog_clk
    PORT
      LAYER met3 ;
        RECT 0.000 6.840 4.000 7.440 ;
    END
  END prog_clk
  PIN right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_
    PORT
      LAYER met2 ;
        RECT 45.170 0.000 45.450 4.000 ;
    END
  END right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_
  PIN right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_
    PORT
      LAYER met2 ;
        RECT 93.470 96.000 93.750 100.000 ;
    END
  END right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_
  PIN right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_
    PORT
      LAYER met2 ;
        RECT 87.030 96.000 87.310 100.000 ;
    END
  END right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_
  PIN right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_
    PORT
      LAYER met2 ;
        RECT 19.410 96.000 19.690 100.000 ;
    END
  END right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_
  PIN right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_
    PORT
      LAYER met2 ;
        RECT 32.290 96.000 32.570 100.000 ;
    END
  END right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_
  PIN right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_
    PORT
      LAYER met2 ;
        RECT 61.270 0.000 61.550 4.000 ;
    END
  END right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_
  PIN right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_
    PORT
      LAYER met3 ;
        RECT 0.000 34.040 4.000 34.640 ;
    END
  END right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_
  PIN right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_
    PORT
      LAYER met3 ;
        RECT 0.000 91.840 4.000 92.440 ;
    END
  END right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_
  PIN right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_
    PORT
      LAYER met3 ;
        RECT 96.000 44.240 100.000 44.840 ;
    END
  END right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_
  PIN vccd1
    PORT
      LAYER met4 ;
        RECT 82.400 10.640 84.000 87.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 60.205 10.640 61.805 87.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 38.010 10.640 39.610 87.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 15.815 10.640 17.415 87.280 ;
    END
  END vccd1
  PIN vssd1
    PORT
      LAYER met4 ;
        RECT 93.495 10.640 95.095 87.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 71.300 10.640 72.900 87.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 49.105 10.640 50.705 87.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 26.910 10.640 28.510 87.280 ;
    END
  END vssd1
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 94.300 87.125 ;
      LAYER met1 ;
        RECT 0.070 8.200 96.070 87.280 ;
      LAYER met2 ;
        RECT 0.100 95.720 6.250 99.125 ;
        RECT 7.090 95.720 12.690 99.125 ;
        RECT 13.530 95.720 19.130 99.125 ;
        RECT 19.970 95.720 25.570 99.125 ;
        RECT 26.410 95.720 32.010 99.125 ;
        RECT 32.850 95.720 38.450 99.125 ;
        RECT 39.290 95.720 44.890 99.125 ;
        RECT 45.730 95.720 54.550 99.125 ;
        RECT 55.390 95.720 60.990 99.125 ;
        RECT 61.830 95.720 67.430 99.125 ;
        RECT 68.270 95.720 73.870 99.125 ;
        RECT 74.710 95.720 80.310 99.125 ;
        RECT 81.150 95.720 86.750 99.125 ;
        RECT 87.590 95.720 93.190 99.125 ;
        RECT 94.030 95.720 96.050 99.125 ;
        RECT 0.100 4.280 96.050 95.720 ;
        RECT 0.650 3.555 6.250 4.280 ;
        RECT 7.090 3.555 12.690 4.280 ;
        RECT 13.530 3.555 19.130 4.280 ;
        RECT 19.970 3.555 25.570 4.280 ;
        RECT 26.410 3.555 32.010 4.280 ;
        RECT 32.850 3.555 38.450 4.280 ;
        RECT 39.290 3.555 44.890 4.280 ;
        RECT 45.730 3.555 54.550 4.280 ;
        RECT 55.390 3.555 60.990 4.280 ;
        RECT 61.830 3.555 67.430 4.280 ;
        RECT 68.270 3.555 73.870 4.280 ;
        RECT 74.710 3.555 80.310 4.280 ;
        RECT 81.150 3.555 86.750 4.280 ;
        RECT 87.590 3.555 93.190 4.280 ;
        RECT 94.030 3.555 96.050 4.280 ;
      LAYER met3 ;
        RECT 4.400 98.240 96.000 99.105 ;
        RECT 4.000 96.240 96.000 98.240 ;
        RECT 4.000 94.840 95.600 96.240 ;
        RECT 4.000 92.840 96.000 94.840 ;
        RECT 4.400 91.440 96.000 92.840 ;
        RECT 4.000 89.440 96.000 91.440 ;
        RECT 4.000 88.040 95.600 89.440 ;
        RECT 4.000 86.040 96.000 88.040 ;
        RECT 4.400 84.640 96.000 86.040 ;
        RECT 4.000 82.640 96.000 84.640 ;
        RECT 4.000 81.240 95.600 82.640 ;
        RECT 4.000 79.240 96.000 81.240 ;
        RECT 4.400 77.840 96.000 79.240 ;
        RECT 4.000 75.840 96.000 77.840 ;
        RECT 4.000 74.440 95.600 75.840 ;
        RECT 4.000 72.440 96.000 74.440 ;
        RECT 4.400 71.040 96.000 72.440 ;
        RECT 4.000 69.040 96.000 71.040 ;
        RECT 4.000 67.640 95.600 69.040 ;
        RECT 4.000 65.640 96.000 67.640 ;
        RECT 4.400 64.240 96.000 65.640 ;
        RECT 4.000 62.240 96.000 64.240 ;
        RECT 4.000 60.840 95.600 62.240 ;
        RECT 4.000 58.840 96.000 60.840 ;
        RECT 4.400 57.440 96.000 58.840 ;
        RECT 4.000 55.440 96.000 57.440 ;
        RECT 4.000 54.040 95.600 55.440 ;
        RECT 4.000 48.640 96.000 54.040 ;
        RECT 4.400 47.240 96.000 48.640 ;
        RECT 4.000 45.240 96.000 47.240 ;
        RECT 4.000 43.840 95.600 45.240 ;
        RECT 4.000 41.840 96.000 43.840 ;
        RECT 4.400 40.440 96.000 41.840 ;
        RECT 4.000 38.440 96.000 40.440 ;
        RECT 4.000 37.040 95.600 38.440 ;
        RECT 4.000 35.040 96.000 37.040 ;
        RECT 4.400 33.640 96.000 35.040 ;
        RECT 4.000 31.640 96.000 33.640 ;
        RECT 4.000 30.240 95.600 31.640 ;
        RECT 4.000 28.240 96.000 30.240 ;
        RECT 4.400 26.840 96.000 28.240 ;
        RECT 4.000 24.840 96.000 26.840 ;
        RECT 4.000 23.440 95.600 24.840 ;
        RECT 4.000 21.440 96.000 23.440 ;
        RECT 4.400 20.040 96.000 21.440 ;
        RECT 4.000 18.040 96.000 20.040 ;
        RECT 4.000 16.640 95.600 18.040 ;
        RECT 4.000 14.640 96.000 16.640 ;
        RECT 4.400 13.240 96.000 14.640 ;
        RECT 4.000 11.240 96.000 13.240 ;
        RECT 4.000 9.840 95.600 11.240 ;
        RECT 4.000 7.840 96.000 9.840 ;
        RECT 4.400 6.440 96.000 7.840 ;
        RECT 4.000 4.440 96.000 6.440 ;
        RECT 4.000 3.575 95.600 4.440 ;
  END
END sb_0__4_
END LIBRARY

