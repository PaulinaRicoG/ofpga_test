VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO cbx_1__4_
  CLASS BLOCK ;
  FOREIGN cbx_1__4_ ;
  ORIGIN 0.000 0.000 ;
  SIZE 100.000 BY 100.000 ;
  PIN bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_
    PORT
      LAYER met3 ;
        RECT 0.000 10.240 4.000 10.840 ;
    END
  END bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_
  PIN bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_
    PORT
      LAYER met3 ;
        RECT 96.000 34.040 100.000 34.640 ;
    END
  END bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_
  PIN bottom_grid_top_width_0_height_0_subtile_0__pin_I0_2_
    PORT
      LAYER met3 ;
        RECT 96.000 3.440 100.000 4.040 ;
    END
  END bottom_grid_top_width_0_height_0_subtile_0__pin_I0_2_
  PIN bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_
    PORT
      LAYER met3 ;
        RECT 0.000 23.840 4.000 24.440 ;
    END
  END bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_
  PIN bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_
    PORT
      LAYER met2 ;
        RECT 41.950 96.000 42.230 100.000 ;
    END
  END bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_
  PIN bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_
    PORT
      LAYER met2 ;
        RECT 19.410 96.000 19.690 100.000 ;
    END
  END bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_
  PIN bottom_grid_top_width_0_height_0_subtile_0__pin_I1_2_
    PORT
      LAYER met2 ;
        RECT 0.090 96.000 0.370 100.000 ;
    END
  END bottom_grid_top_width_0_height_0_subtile_0__pin_I1_2_
  PIN bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_
    PORT
      LAYER met3 ;
        RECT 0.000 64.640 4.000 65.240 ;
    END
  END bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_
  PIN bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_
    PORT
      LAYER met3 ;
        RECT 96.000 68.040 100.000 68.640 ;
    END
  END bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_
  PIN bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_
    PORT
      LAYER met3 ;
        RECT 96.000 17.040 100.000 17.640 ;
    END
  END bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_
  PIN bottom_grid_top_width_0_height_0_subtile_0__pin_I2_2_
    PORT
      LAYER met2 ;
        RECT 22.630 0.000 22.910 4.000 ;
    END
  END bottom_grid_top_width_0_height_0_subtile_0__pin_I2_2_
  PIN bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_
    PORT
      LAYER met2 ;
        RECT 35.510 96.000 35.790 100.000 ;
    END
  END bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_
  PIN bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_
    PORT
      LAYER met2 ;
        RECT 67.710 96.000 67.990 100.000 ;
    END
  END bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_
  PIN bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_
    PORT
      LAYER met2 ;
        RECT 61.270 0.000 61.550 4.000 ;
    END
  END bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_
  PIN bottom_grid_top_width_0_height_0_subtile_0__pin_I3_2_
    PORT
      LAYER met2 ;
        RECT 3.310 0.000 3.590 4.000 ;
    END
  END bottom_grid_top_width_0_height_0_subtile_0__pin_I3_2_
  PIN bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_
    PORT
      LAYER met3 ;
        RECT 96.000 54.440 100.000 55.040 ;
    END
  END bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_
  PIN ccff_head
    PORT
      LAYER met3 ;
        RECT 96.000 30.640 100.000 31.240 ;
    END
  END ccff_head
  PIN ccff_tail
    PORT
      LAYER met2 ;
        RECT 54.830 96.000 55.110 100.000 ;
    END
  END ccff_tail
  PIN chanx_left_in[0]
    PORT
      LAYER met3 ;
        RECT 96.000 88.440 100.000 89.040 ;
    END
  END chanx_left_in[0]
  PIN chanx_left_in[10]
    PORT
      LAYER met3 ;
        RECT 0.000 74.840 4.000 75.440 ;
    END
  END chanx_left_in[10]
  PIN chanx_left_in[1]
    PORT
      LAYER met3 ;
        RECT 96.000 61.240 100.000 61.840 ;
    END
  END chanx_left_in[1]
  PIN chanx_left_in[2]
    PORT
      LAYER met3 ;
        RECT 0.000 81.640 4.000 82.240 ;
    END
  END chanx_left_in[2]
  PIN chanx_left_in[3]
    PORT
      LAYER met3 ;
        RECT 96.000 95.240 100.000 95.840 ;
    END
  END chanx_left_in[3]
  PIN chanx_left_in[4]
    PORT
      LAYER met2 ;
        RECT 83.810 0.000 84.090 4.000 ;
    END
  END chanx_left_in[4]
  PIN chanx_left_in[5]
    PORT
      LAYER met2 ;
        RECT 77.370 0.000 77.650 4.000 ;
    END
  END chanx_left_in[5]
  PIN chanx_left_in[6]
    PORT
      LAYER met2 ;
        RECT 41.950 0.000 42.230 4.000 ;
    END
  END chanx_left_in[6]
  PIN chanx_left_in[7]
    PORT
      LAYER met2 ;
        RECT 6.530 96.000 6.810 100.000 ;
    END
  END chanx_left_in[7]
  PIN chanx_left_in[8]
    PORT
      LAYER met2 ;
        RECT 70.930 0.000 71.210 4.000 ;
    END
  END chanx_left_in[8]
  PIN chanx_left_in[9]
    PORT
      LAYER met2 ;
        RECT 61.270 96.000 61.550 100.000 ;
    END
  END chanx_left_in[9]
  PIN chanx_left_out[0]
    PORT
      LAYER met2 ;
        RECT 90.250 0.000 90.530 4.000 ;
    END
  END chanx_left_out[0]
  PIN chanx_left_out[10]
    PORT
      LAYER met3 ;
        RECT 96.000 10.240 100.000 10.840 ;
    END
  END chanx_left_out[10]
  PIN chanx_left_out[1]
    PORT
      LAYER met2 ;
        RECT 54.830 0.000 55.110 4.000 ;
    END
  END chanx_left_out[1]
  PIN chanx_left_out[2]
    PORT
      LAYER met3 ;
        RECT 96.000 23.840 100.000 24.440 ;
    END
  END chanx_left_out[2]
  PIN chanx_left_out[3]
    PORT
      LAYER met2 ;
        RECT 80.590 96.000 80.870 100.000 ;
    END
  END chanx_left_out[3]
  PIN chanx_left_out[4]
    PORT
      LAYER met3 ;
        RECT 0.000 51.040 4.000 51.640 ;
    END
  END chanx_left_out[4]
  PIN chanx_left_out[5]
    PORT
      LAYER met3 ;
        RECT 0.000 17.040 4.000 17.640 ;
    END
  END chanx_left_out[5]
  PIN chanx_left_out[6]
    PORT
      LAYER met3 ;
        RECT 0.000 95.240 4.000 95.840 ;
    END
  END chanx_left_out[6]
  PIN chanx_left_out[7]
    PORT
      LAYER met3 ;
        RECT 0.000 68.040 4.000 68.640 ;
    END
  END chanx_left_out[7]
  PIN chanx_left_out[8]
    PORT
      LAYER met2 ;
        RECT 74.150 96.000 74.430 100.000 ;
    END
  END chanx_left_out[8]
  PIN chanx_left_out[9]
    PORT
      LAYER met2 ;
        RECT 93.470 96.000 93.750 100.000 ;
    END
  END chanx_left_out[9]
  PIN chanx_right_in[0]
    PORT
      LAYER met2 ;
        RECT 25.850 96.000 26.130 100.000 ;
    END
  END chanx_right_in[0]
  PIN chanx_right_in[10]
    PORT
      LAYER met2 ;
        RECT 48.390 96.000 48.670 100.000 ;
    END
  END chanx_right_in[10]
  PIN chanx_right_in[1]
    PORT
      LAYER met2 ;
        RECT 9.750 0.000 10.030 4.000 ;
    END
  END chanx_right_in[1]
  PIN chanx_right_in[2]
    PORT
      LAYER met2 ;
        RECT 0.090 0.000 0.370 4.000 ;
    END
  END chanx_right_in[2]
  PIN chanx_right_in[3]
    PORT
      LAYER met3 ;
        RECT 96.000 81.640 100.000 82.240 ;
    END
  END chanx_right_in[3]
  PIN chanx_right_in[4]
    PORT
      LAYER met2 ;
        RECT 96.690 96.000 96.970 100.000 ;
    END
  END chanx_right_in[4]
  PIN chanx_right_in[5]
    PORT
      LAYER met2 ;
        RECT 35.510 0.000 35.790 4.000 ;
    END
  END chanx_right_in[5]
  PIN chanx_right_in[6]
    PORT
      LAYER met3 ;
        RECT 96.000 74.840 100.000 75.440 ;
    END
  END chanx_right_in[6]
  PIN chanx_right_in[7]
    PORT
      LAYER met2 ;
        RECT 96.690 0.000 96.970 4.000 ;
    END
  END chanx_right_in[7]
  PIN chanx_right_in[8]
    PORT
      LAYER met3 ;
        RECT 0.000 30.640 4.000 31.240 ;
    END
  END chanx_right_in[8]
  PIN chanx_right_in[9]
    PORT
      LAYER met3 ;
        RECT 0.000 3.440 4.000 4.040 ;
    END
  END chanx_right_in[9]
  PIN chanx_right_out[0]
    PORT
      LAYER met2 ;
        RECT 16.190 0.000 16.470 4.000 ;
    END
  END chanx_right_out[0]
  PIN chanx_right_out[10]
    PORT
      LAYER met2 ;
        RECT 29.070 0.000 29.350 4.000 ;
    END
  END chanx_right_out[10]
  PIN chanx_right_out[1]
    PORT
      LAYER met3 ;
        RECT 0.000 57.840 4.000 58.440 ;
    END
  END chanx_right_out[1]
  PIN chanx_right_out[2]
    PORT
      LAYER met3 ;
        RECT 96.000 47.640 100.000 48.240 ;
    END
  END chanx_right_out[2]
  PIN chanx_right_out[3]
    PORT
      LAYER met2 ;
        RECT 48.390 0.000 48.670 4.000 ;
    END
  END chanx_right_out[3]
  PIN chanx_right_out[4]
    PORT
      LAYER met3 ;
        RECT 0.000 44.240 4.000 44.840 ;
    END
  END chanx_right_out[4]
  PIN chanx_right_out[5]
    PORT
      LAYER met2 ;
        RECT 87.030 96.000 87.310 100.000 ;
    END
  END chanx_right_out[5]
  PIN chanx_right_out[6]
    PORT
      LAYER met2 ;
        RECT 12.970 96.000 13.250 100.000 ;
    END
  END chanx_right_out[6]
  PIN chanx_right_out[7]
    PORT
      LAYER met2 ;
        RECT 32.290 96.000 32.570 100.000 ;
    END
  END chanx_right_out[7]
  PIN chanx_right_out[8]
    PORT
      LAYER met2 ;
        RECT 64.490 0.000 64.770 4.000 ;
    END
  END chanx_right_out[8]
  PIN chanx_right_out[9]
    PORT
      LAYER met3 ;
        RECT 0.000 37.440 4.000 38.040 ;
    END
  END chanx_right_out[9]
  PIN prog_clk
    PORT
      LAYER met3 ;
        RECT 0.000 88.440 4.000 89.040 ;
    END
  END prog_clk
  PIN top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_
    PORT
      LAYER met3 ;
        RECT 96.000 40.840 100.000 41.440 ;
    END
  END top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_
  PIN vccd1
    PORT
      LAYER met4 ;
        RECT 82.400 10.640 84.000 87.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 60.205 10.640 61.805 87.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 38.010 10.640 39.610 87.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 15.815 10.640 17.415 87.280 ;
    END
  END vccd1
  PIN vssd1
    PORT
      LAYER met4 ;
        RECT 93.495 10.640 95.095 87.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 71.300 10.640 72.900 87.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 49.105 10.640 50.705 87.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 26.910 10.640 28.510 87.280 ;
    END
  END vssd1
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 94.300 87.125 ;
      LAYER met1 ;
        RECT 0.070 10.640 96.990 89.380 ;
      LAYER met2 ;
        RECT 0.650 95.720 6.250 96.290 ;
        RECT 7.090 95.720 12.690 96.290 ;
        RECT 13.530 95.720 19.130 96.290 ;
        RECT 19.970 95.720 25.570 96.290 ;
        RECT 26.410 95.720 32.010 96.290 ;
        RECT 32.850 95.720 35.230 96.290 ;
        RECT 36.070 95.720 41.670 96.290 ;
        RECT 42.510 95.720 48.110 96.290 ;
        RECT 48.950 95.720 54.550 96.290 ;
        RECT 55.390 95.720 60.990 96.290 ;
        RECT 61.830 95.720 67.430 96.290 ;
        RECT 68.270 95.720 73.870 96.290 ;
        RECT 74.710 95.720 80.310 96.290 ;
        RECT 81.150 95.720 86.750 96.290 ;
        RECT 87.590 95.720 93.190 96.290 ;
        RECT 94.030 95.720 96.410 96.290 ;
        RECT 0.100 4.280 96.960 95.720 ;
        RECT 0.650 3.555 3.030 4.280 ;
        RECT 3.870 3.555 9.470 4.280 ;
        RECT 10.310 3.555 15.910 4.280 ;
        RECT 16.750 3.555 22.350 4.280 ;
        RECT 23.190 3.555 28.790 4.280 ;
        RECT 29.630 3.555 35.230 4.280 ;
        RECT 36.070 3.555 41.670 4.280 ;
        RECT 42.510 3.555 48.110 4.280 ;
        RECT 48.950 3.555 54.550 4.280 ;
        RECT 55.390 3.555 60.990 4.280 ;
        RECT 61.830 3.555 64.210 4.280 ;
        RECT 65.050 3.555 70.650 4.280 ;
        RECT 71.490 3.555 77.090 4.280 ;
        RECT 77.930 3.555 83.530 4.280 ;
        RECT 84.370 3.555 89.970 4.280 ;
        RECT 90.810 3.555 96.410 4.280 ;
      LAYER met3 ;
        RECT 4.400 94.840 95.600 95.705 ;
        RECT 4.000 89.440 96.000 94.840 ;
        RECT 4.400 88.040 95.600 89.440 ;
        RECT 4.000 82.640 96.000 88.040 ;
        RECT 4.400 81.240 95.600 82.640 ;
        RECT 4.000 75.840 96.000 81.240 ;
        RECT 4.400 74.440 95.600 75.840 ;
        RECT 4.000 69.040 96.000 74.440 ;
        RECT 4.400 67.640 95.600 69.040 ;
        RECT 4.000 65.640 96.000 67.640 ;
        RECT 4.400 64.240 96.000 65.640 ;
        RECT 4.000 62.240 96.000 64.240 ;
        RECT 4.000 60.840 95.600 62.240 ;
        RECT 4.000 58.840 96.000 60.840 ;
        RECT 4.400 57.440 96.000 58.840 ;
        RECT 4.000 55.440 96.000 57.440 ;
        RECT 4.000 54.040 95.600 55.440 ;
        RECT 4.000 52.040 96.000 54.040 ;
        RECT 4.400 50.640 96.000 52.040 ;
        RECT 4.000 48.640 96.000 50.640 ;
        RECT 4.000 47.240 95.600 48.640 ;
        RECT 4.000 45.240 96.000 47.240 ;
        RECT 4.400 43.840 96.000 45.240 ;
        RECT 4.000 41.840 96.000 43.840 ;
        RECT 4.000 40.440 95.600 41.840 ;
        RECT 4.000 38.440 96.000 40.440 ;
        RECT 4.400 37.040 96.000 38.440 ;
        RECT 4.000 35.040 96.000 37.040 ;
        RECT 4.000 33.640 95.600 35.040 ;
        RECT 4.000 31.640 96.000 33.640 ;
        RECT 4.400 30.240 95.600 31.640 ;
        RECT 4.000 24.840 96.000 30.240 ;
        RECT 4.400 23.440 95.600 24.840 ;
        RECT 4.000 18.040 96.000 23.440 ;
        RECT 4.400 16.640 95.600 18.040 ;
        RECT 4.000 11.240 96.000 16.640 ;
        RECT 4.400 9.840 95.600 11.240 ;
        RECT 4.000 4.440 96.000 9.840 ;
        RECT 4.400 3.575 95.600 4.440 ;
      LAYER met4 ;
        RECT 17.775 87.680 76.065 89.585 ;
        RECT 17.815 36.895 26.510 87.680 ;
        RECT 28.910 36.895 37.610 87.680 ;
        RECT 40.010 36.895 48.705 87.680 ;
        RECT 51.105 36.895 59.805 87.680 ;
        RECT 62.205 36.895 70.900 87.680 ;
        RECT 73.300 36.895 76.065 87.680 ;
  END
END cbx_1__4_
END LIBRARY

