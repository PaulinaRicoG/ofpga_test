VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO grid_clb
  CLASS BLOCK ;
  FOREIGN grid_clb ;
  ORIGIN 0.000 0.000 ;
  SIZE 110.000 BY 110.000 ;
  PIN Test_en
    PORT
      LAYER met3 ;
        RECT 106.000 88.440 110.000 89.040 ;
    END
  END Test_en
  PIN bottom_width_0_height_0_subtile_0__pin_regout_0_
    PORT
      LAYER met3 ;
        RECT 106.000 57.840 110.000 58.440 ;
    END
  END bottom_width_0_height_0_subtile_0__pin_regout_0_
  PIN bottom_width_0_height_0_subtile_0__pin_scout_0_
    PORT
      LAYER met2 ;
        RECT 64.490 0.000 64.770 4.000 ;
    END
  END bottom_width_0_height_0_subtile_0__pin_scout_0_
  PIN ccff_head
    PORT
      LAYER met3 ;
        RECT 0.000 13.640 4.000 14.240 ;
    END
  END ccff_head
  PIN ccff_tail
    PORT
      LAYER met2 ;
        RECT 9.750 106.000 10.030 110.000 ;
    END
  END ccff_tail
  PIN clk
    PORT
      LAYER met3 ;
        RECT 106.000 27.240 110.000 27.840 ;
    END
  END clk
  PIN left_width_0_height_0_subtile_0__pin_clk_0_
    PORT
      LAYER met3 ;
        RECT 106.000 95.240 110.000 95.840 ;
    END
  END left_width_0_height_0_subtile_0__pin_clk_0_
  PIN prog_clk
    PORT
      LAYER met2 ;
        RECT 6.530 0.000 6.810 4.000 ;
    END
  END prog_clk
  PIN reset
    PORT
      LAYER met3 ;
        RECT 106.000 34.040 110.000 34.640 ;
    END
  END reset
  PIN right_width_0_height_0_subtile_0__pin_I4_0_
    PORT
      LAYER met3 ;
        RECT 106.000 17.040 110.000 17.640 ;
    END
  END right_width_0_height_0_subtile_0__pin_I4_0_
  PIN right_width_0_height_0_subtile_0__pin_I4_1_
    PORT
      LAYER met2 ;
        RECT 61.270 106.000 61.550 110.000 ;
    END
  END right_width_0_height_0_subtile_0__pin_I4_1_
  PIN right_width_0_height_0_subtile_0__pin_I4_2_
    PORT
      LAYER met3 ;
        RECT 106.000 71.440 110.000 72.040 ;
    END
  END right_width_0_height_0_subtile_0__pin_I4_2_
  PIN right_width_0_height_0_subtile_0__pin_I4i_0_
    PORT
      LAYER met2 ;
        RECT 19.410 0.000 19.690 4.000 ;
    END
  END right_width_0_height_0_subtile_0__pin_I4i_0_
  PIN right_width_0_height_0_subtile_0__pin_I5_0_
    PORT
      LAYER met2 ;
        RECT 74.150 106.000 74.430 110.000 ;
    END
  END right_width_0_height_0_subtile_0__pin_I5_0_
  PIN right_width_0_height_0_subtile_0__pin_I5_1_
    PORT
      LAYER met2 ;
        RECT 99.910 0.000 100.190 4.000 ;
    END
  END right_width_0_height_0_subtile_0__pin_I5_1_
  PIN right_width_0_height_0_subtile_0__pin_I5_2_
    PORT
      LAYER met3 ;
        RECT 0.000 91.840 4.000 92.440 ;
    END
  END right_width_0_height_0_subtile_0__pin_I5_2_
  PIN right_width_0_height_0_subtile_0__pin_I5i_0_
    PORT
      LAYER met3 ;
        RECT 0.000 74.840 4.000 75.440 ;
    END
  END right_width_0_height_0_subtile_0__pin_I5i_0_
  PIN right_width_0_height_0_subtile_0__pin_I6_0_
    PORT
      LAYER met2 ;
        RECT 51.610 106.000 51.890 110.000 ;
    END
  END right_width_0_height_0_subtile_0__pin_I6_0_
  PIN right_width_0_height_0_subtile_0__pin_I6_1_
    PORT
      LAYER met2 ;
        RECT 90.250 106.000 90.530 110.000 ;
    END
  END right_width_0_height_0_subtile_0__pin_I6_1_
  PIN right_width_0_height_0_subtile_0__pin_I6_2_
    PORT
      LAYER met2 ;
        RECT 87.030 0.000 87.310 4.000 ;
    END
  END right_width_0_height_0_subtile_0__pin_I6_2_
  PIN right_width_0_height_0_subtile_0__pin_I6i_0_
    PORT
      LAYER met2 ;
        RECT 77.370 0.000 77.650 4.000 ;
    END
  END right_width_0_height_0_subtile_0__pin_I6i_0_
  PIN right_width_0_height_0_subtile_0__pin_I7_0_
    PORT
      LAYER met3 ;
        RECT 0.000 44.240 4.000 44.840 ;
    END
  END right_width_0_height_0_subtile_0__pin_I7_0_
  PIN right_width_0_height_0_subtile_0__pin_I7_1_
    PORT
      LAYER met3 ;
        RECT 106.000 64.640 110.000 65.240 ;
    END
  END right_width_0_height_0_subtile_0__pin_I7_1_
  PIN right_width_0_height_0_subtile_0__pin_I7_2_
    PORT
      LAYER met3 ;
        RECT 0.000 30.640 4.000 31.240 ;
    END
  END right_width_0_height_0_subtile_0__pin_I7_2_
  PIN right_width_0_height_0_subtile_0__pin_I7i_0_
    PORT
      LAYER met2 ;
        RECT 80.590 106.000 80.870 110.000 ;
    END
  END right_width_0_height_0_subtile_0__pin_I7i_0_
  PIN right_width_0_height_0_subtile_0__pin_O_10_
    PORT
      LAYER met2 ;
        RECT 93.470 0.000 93.750 4.000 ;
    END
  END right_width_0_height_0_subtile_0__pin_O_10_
  PIN right_width_0_height_0_subtile_0__pin_O_11_
    PORT
      LAYER met3 ;
        RECT 106.000 3.440 110.000 4.040 ;
    END
  END right_width_0_height_0_subtile_0__pin_O_11_
  PIN right_width_0_height_0_subtile_0__pin_O_12_
    PORT
      LAYER met3 ;
        RECT 0.000 68.040 4.000 68.640 ;
    END
  END right_width_0_height_0_subtile_0__pin_O_12_
  PIN right_width_0_height_0_subtile_0__pin_O_13_
    PORT
      LAYER met3 ;
        RECT 106.000 10.240 110.000 10.840 ;
    END
  END right_width_0_height_0_subtile_0__pin_O_13_
  PIN right_width_0_height_0_subtile_0__pin_O_14_
    PORT
      LAYER met3 ;
        RECT 0.000 61.240 4.000 61.840 ;
    END
  END right_width_0_height_0_subtile_0__pin_O_14_
  PIN right_width_0_height_0_subtile_0__pin_O_15_
    PORT
      LAYER met2 ;
        RECT 109.570 106.000 109.850 110.000 ;
    END
  END right_width_0_height_0_subtile_0__pin_O_15_
  PIN right_width_0_height_0_subtile_0__pin_O_8_
    PORT
      LAYER met2 ;
        RECT 35.510 0.000 35.790 4.000 ;
    END
  END right_width_0_height_0_subtile_0__pin_O_8_
  PIN right_width_0_height_0_subtile_0__pin_O_9_
    PORT
      LAYER met2 ;
        RECT 0.090 106.000 0.370 110.000 ;
    END
  END right_width_0_height_0_subtile_0__pin_O_9_
  PIN set
    PORT
      LAYER met3 ;
        RECT 0.000 81.640 4.000 82.240 ;
    END
  END set
  PIN top_width_0_height_0_subtile_0__pin_I0_0_
    PORT
      LAYER met3 ;
        RECT 0.000 51.040 4.000 51.640 ;
    END
  END top_width_0_height_0_subtile_0__pin_I0_0_
  PIN top_width_0_height_0_subtile_0__pin_I0_1_
    PORT
      LAYER met2 ;
        RECT 32.290 106.000 32.570 110.000 ;
    END
  END top_width_0_height_0_subtile_0__pin_I0_1_
  PIN top_width_0_height_0_subtile_0__pin_I0_2_
    PORT
      LAYER met3 ;
        RECT 0.000 20.440 4.000 21.040 ;
    END
  END top_width_0_height_0_subtile_0__pin_I0_2_
  PIN top_width_0_height_0_subtile_0__pin_I0i_0_
    PORT
      LAYER met2 ;
        RECT 67.710 106.000 67.990 110.000 ;
    END
  END top_width_0_height_0_subtile_0__pin_I0i_0_
  PIN top_width_0_height_0_subtile_0__pin_I1_0_
    PORT
      LAYER met3 ;
        RECT 0.000 98.640 4.000 99.240 ;
    END
  END top_width_0_height_0_subtile_0__pin_I1_0_
  PIN top_width_0_height_0_subtile_0__pin_I1_1_
    PORT
      LAYER met2 ;
        RECT 0.090 0.000 0.370 4.000 ;
    END
  END top_width_0_height_0_subtile_0__pin_I1_1_
  PIN top_width_0_height_0_subtile_0__pin_I1_2_
    PORT
      LAYER met2 ;
        RECT 16.190 106.000 16.470 110.000 ;
    END
  END top_width_0_height_0_subtile_0__pin_I1_2_
  PIN top_width_0_height_0_subtile_0__pin_I1i_0_
    PORT
      LAYER met3 ;
        RECT 106.000 102.040 110.000 102.640 ;
    END
  END top_width_0_height_0_subtile_0__pin_I1i_0_
  PIN top_width_0_height_0_subtile_0__pin_I2_0_
    PORT
      LAYER met2 ;
        RECT 41.950 0.000 42.230 4.000 ;
    END
  END top_width_0_height_0_subtile_0__pin_I2_0_
  PIN top_width_0_height_0_subtile_0__pin_I2_1_
    PORT
      LAYER met3 ;
        RECT 106.000 78.240 110.000 78.840 ;
    END
  END top_width_0_height_0_subtile_0__pin_I2_1_
  PIN top_width_0_height_0_subtile_0__pin_I2_2_
    PORT
      LAYER met2 ;
        RECT 109.570 0.000 109.850 4.000 ;
    END
  END top_width_0_height_0_subtile_0__pin_I2_2_
  PIN top_width_0_height_0_subtile_0__pin_I2i_0_
    PORT
      LAYER met2 ;
        RECT 45.170 106.000 45.450 110.000 ;
    END
  END top_width_0_height_0_subtile_0__pin_I2i_0_
  PIN top_width_0_height_0_subtile_0__pin_I3_0_
    PORT
      LAYER met3 ;
        RECT 106.000 40.840 110.000 41.440 ;
    END
  END top_width_0_height_0_subtile_0__pin_I3_0_
  PIN top_width_0_height_0_subtile_0__pin_I3_1_
    PORT
      LAYER met2 ;
        RECT 12.970 0.000 13.250 4.000 ;
    END
  END top_width_0_height_0_subtile_0__pin_I3_1_
  PIN top_width_0_height_0_subtile_0__pin_I3_2_
    PORT
      LAYER met2 ;
        RECT 29.070 0.000 29.350 4.000 ;
    END
  END top_width_0_height_0_subtile_0__pin_I3_2_
  PIN top_width_0_height_0_subtile_0__pin_I3i_0_
    PORT
      LAYER met2 ;
        RECT 48.390 0.000 48.670 4.000 ;
    END
  END top_width_0_height_0_subtile_0__pin_I3i_0_
  PIN top_width_0_height_0_subtile_0__pin_O_0_
    PORT
      LAYER met3 ;
        RECT 0.000 6.840 4.000 7.440 ;
    END
  END top_width_0_height_0_subtile_0__pin_O_0_
  PIN top_width_0_height_0_subtile_0__pin_O_1_
    PORT
      LAYER met2 ;
        RECT 58.050 0.000 58.330 4.000 ;
    END
  END top_width_0_height_0_subtile_0__pin_O_1_
  PIN top_width_0_height_0_subtile_0__pin_O_2_
    PORT
      LAYER met2 ;
        RECT 103.130 106.000 103.410 110.000 ;
    END
  END top_width_0_height_0_subtile_0__pin_O_2_
  PIN top_width_0_height_0_subtile_0__pin_O_3_
    PORT
      LAYER met2 ;
        RECT 96.690 106.000 96.970 110.000 ;
    END
  END top_width_0_height_0_subtile_0__pin_O_3_
  PIN top_width_0_height_0_subtile_0__pin_O_4_
    PORT
      LAYER met2 ;
        RECT 22.630 106.000 22.910 110.000 ;
    END
  END top_width_0_height_0_subtile_0__pin_O_4_
  PIN top_width_0_height_0_subtile_0__pin_O_5_
    PORT
      LAYER met2 ;
        RECT 38.730 106.000 39.010 110.000 ;
    END
  END top_width_0_height_0_subtile_0__pin_O_5_
  PIN top_width_0_height_0_subtile_0__pin_O_6_
    PORT
      LAYER met2 ;
        RECT 70.930 0.000 71.210 4.000 ;
    END
  END top_width_0_height_0_subtile_0__pin_O_6_
  PIN top_width_0_height_0_subtile_0__pin_O_7_
    PORT
      LAYER met3 ;
        RECT 0.000 37.440 4.000 38.040 ;
    END
  END top_width_0_height_0_subtile_0__pin_O_7_
  PIN top_width_0_height_0_subtile_0__pin_regin_0_
    PORT
      LAYER met3 ;
        RECT 0.000 105.440 4.000 106.040 ;
    END
  END top_width_0_height_0_subtile_0__pin_regin_0_
  PIN top_width_0_height_0_subtile_0__pin_scin_0_
    PORT
      LAYER met3 ;
        RECT 106.000 47.640 110.000 48.240 ;
    END
  END top_width_0_height_0_subtile_0__pin_scin_0_
  PIN vccd1
    PORT
      LAYER met4 ;
        RECT 91.255 10.640 92.855 98.160 ;
    END
    PORT
      LAYER met4 ;
        RECT 66.530 10.640 68.130 98.160 ;
    END
    PORT
      LAYER met4 ;
        RECT 41.805 10.640 43.405 98.160 ;
    END
    PORT
      LAYER met4 ;
        RECT 17.080 10.640 18.680 98.160 ;
    END
  END vccd1
  PIN vssd1
    PORT
      LAYER met4 ;
        RECT 103.615 10.640 105.215 98.160 ;
    END
    PORT
      LAYER met4 ;
        RECT 78.890 10.640 80.490 98.160 ;
    END
    PORT
      LAYER met4 ;
        RECT 54.165 10.640 55.765 98.160 ;
    END
    PORT
      LAYER met4 ;
        RECT 29.440 10.640 31.040 98.160 ;
    END
  END vssd1
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 104.420 98.005 ;
      LAYER met1 ;
        RECT 0.070 9.220 109.870 99.240 ;
      LAYER met2 ;
        RECT 0.650 105.720 9.470 106.490 ;
        RECT 10.310 105.720 15.910 106.490 ;
        RECT 16.750 105.720 22.350 106.490 ;
        RECT 23.190 105.720 32.010 106.490 ;
        RECT 32.850 105.720 38.450 106.490 ;
        RECT 39.290 105.720 44.890 106.490 ;
        RECT 45.730 105.720 51.330 106.490 ;
        RECT 52.170 105.720 60.990 106.490 ;
        RECT 61.830 105.720 67.430 106.490 ;
        RECT 68.270 105.720 73.870 106.490 ;
        RECT 74.710 105.720 80.310 106.490 ;
        RECT 81.150 105.720 89.970 106.490 ;
        RECT 90.810 105.720 96.410 106.490 ;
        RECT 97.250 105.720 102.850 106.490 ;
        RECT 103.690 105.720 109.290 106.490 ;
        RECT 0.100 4.280 109.840 105.720 ;
        RECT 0.650 3.555 6.250 4.280 ;
        RECT 7.090 3.555 12.690 4.280 ;
        RECT 13.530 3.555 19.130 4.280 ;
        RECT 19.970 3.555 28.790 4.280 ;
        RECT 29.630 3.555 35.230 4.280 ;
        RECT 36.070 3.555 41.670 4.280 ;
        RECT 42.510 3.555 48.110 4.280 ;
        RECT 48.950 3.555 57.770 4.280 ;
        RECT 58.610 3.555 64.210 4.280 ;
        RECT 65.050 3.555 70.650 4.280 ;
        RECT 71.490 3.555 77.090 4.280 ;
        RECT 77.930 3.555 86.750 4.280 ;
        RECT 87.590 3.555 93.190 4.280 ;
        RECT 94.030 3.555 99.630 4.280 ;
        RECT 100.470 3.555 109.290 4.280 ;
      LAYER met3 ;
        RECT 4.400 105.040 106.410 105.905 ;
        RECT 4.000 103.040 106.410 105.040 ;
        RECT 4.000 101.640 105.600 103.040 ;
        RECT 4.000 99.640 106.410 101.640 ;
        RECT 4.400 98.240 106.410 99.640 ;
        RECT 4.000 96.240 106.410 98.240 ;
        RECT 4.000 94.840 105.600 96.240 ;
        RECT 4.000 92.840 106.410 94.840 ;
        RECT 4.400 91.440 106.410 92.840 ;
        RECT 4.000 89.440 106.410 91.440 ;
        RECT 4.000 88.040 105.600 89.440 ;
        RECT 4.000 82.640 106.410 88.040 ;
        RECT 4.400 81.240 106.410 82.640 ;
        RECT 4.000 79.240 106.410 81.240 ;
        RECT 4.000 77.840 105.600 79.240 ;
        RECT 4.000 75.840 106.410 77.840 ;
        RECT 4.400 74.440 106.410 75.840 ;
        RECT 4.000 72.440 106.410 74.440 ;
        RECT 4.000 71.040 105.600 72.440 ;
        RECT 4.000 69.040 106.410 71.040 ;
        RECT 4.400 67.640 106.410 69.040 ;
        RECT 4.000 65.640 106.410 67.640 ;
        RECT 4.000 64.240 105.600 65.640 ;
        RECT 4.000 62.240 106.410 64.240 ;
        RECT 4.400 60.840 106.410 62.240 ;
        RECT 4.000 58.840 106.410 60.840 ;
        RECT 4.000 57.440 105.600 58.840 ;
        RECT 4.000 52.040 106.410 57.440 ;
        RECT 4.400 50.640 106.410 52.040 ;
        RECT 4.000 48.640 106.410 50.640 ;
        RECT 4.000 47.240 105.600 48.640 ;
        RECT 4.000 45.240 106.410 47.240 ;
        RECT 4.400 43.840 106.410 45.240 ;
        RECT 4.000 41.840 106.410 43.840 ;
        RECT 4.000 40.440 105.600 41.840 ;
        RECT 4.000 38.440 106.410 40.440 ;
        RECT 4.400 37.040 106.410 38.440 ;
        RECT 4.000 35.040 106.410 37.040 ;
        RECT 4.000 33.640 105.600 35.040 ;
        RECT 4.000 31.640 106.410 33.640 ;
        RECT 4.400 30.240 106.410 31.640 ;
        RECT 4.000 28.240 106.410 30.240 ;
        RECT 4.000 26.840 105.600 28.240 ;
        RECT 4.000 21.440 106.410 26.840 ;
        RECT 4.400 20.040 106.410 21.440 ;
        RECT 4.000 18.040 106.410 20.040 ;
        RECT 4.000 16.640 105.600 18.040 ;
        RECT 4.000 14.640 106.410 16.640 ;
        RECT 4.400 13.240 106.410 14.640 ;
        RECT 4.000 11.240 106.410 13.240 ;
        RECT 4.000 9.840 105.600 11.240 ;
        RECT 4.000 7.840 106.410 9.840 ;
        RECT 4.400 6.440 106.410 7.840 ;
        RECT 4.000 4.440 106.410 6.440 ;
        RECT 4.000 3.575 105.600 4.440 ;
      LAYER met4 ;
        RECT 75.735 17.175 78.490 86.865 ;
        RECT 80.890 17.175 90.785 86.865 ;
  END
END grid_clb
END LIBRARY

