VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO cby_0__1_
  CLASS BLOCK ;
  FOREIGN cby_0__1_ ;
  ORIGIN 0.000 0.000 ;
  SIZE 100.000 BY 100.000 ;
  PIN ccff_head
    PORT
      LAYER met2 ;
        RECT 6.530 96.000 6.810 100.000 ;
    END
  END ccff_head
  PIN ccff_tail
    PORT
      LAYER met3 ;
        RECT 0.000 30.640 4.000 31.240 ;
    END
  END ccff_tail
  PIN chany_bottom_in[0]
    PORT
      LAYER met3 ;
        RECT 96.000 88.440 100.000 89.040 ;
    END
  END chany_bottom_in[0]
  PIN chany_bottom_in[10]
    PORT
      LAYER met3 ;
        RECT 96.000 10.240 100.000 10.840 ;
    END
  END chany_bottom_in[10]
  PIN chany_bottom_in[1]
    PORT
      LAYER met2 ;
        RECT 77.370 96.000 77.650 100.000 ;
    END
  END chany_bottom_in[1]
  PIN chany_bottom_in[2]
    PORT
      LAYER met3 ;
        RECT 0.000 13.640 4.000 14.240 ;
    END
  END chany_bottom_in[2]
  PIN chany_bottom_in[3]
    PORT
      LAYER met3 ;
        RECT 0.000 81.640 4.000 82.240 ;
    END
  END chany_bottom_in[3]
  PIN chany_bottom_in[4]
    PORT
      LAYER met2 ;
        RECT 77.370 0.000 77.650 4.000 ;
    END
  END chany_bottom_in[4]
  PIN chany_bottom_in[5]
    PORT
      LAYER met3 ;
        RECT 96.000 20.440 100.000 21.040 ;
    END
  END chany_bottom_in[5]
  PIN chany_bottom_in[6]
    PORT
      LAYER met2 ;
        RECT 93.470 0.000 93.750 4.000 ;
    END
  END chany_bottom_in[6]
  PIN chany_bottom_in[7]
    PORT
      LAYER met3 ;
        RECT 0.000 64.640 4.000 65.240 ;
    END
  END chany_bottom_in[7]
  PIN chany_bottom_in[8]
    PORT
      LAYER met3 ;
        RECT 96.000 3.440 100.000 4.040 ;
    END
  END chany_bottom_in[8]
  PIN chany_bottom_in[9]
    PORT
      LAYER met2 ;
        RECT 12.970 96.000 13.250 100.000 ;
    END
  END chany_bottom_in[9]
  PIN chany_bottom_out[0]
    PORT
      LAYER met3 ;
        RECT 0.000 47.640 4.000 48.240 ;
    END
  END chany_bottom_out[0]
  PIN chany_bottom_out[10]
    PORT
      LAYER met2 ;
        RECT 54.830 0.000 55.110 4.000 ;
    END
  END chany_bottom_out[10]
  PIN chany_bottom_out[1]
    PORT
      LAYER met2 ;
        RECT 70.930 0.000 71.210 4.000 ;
    END
  END chany_bottom_out[1]
  PIN chany_bottom_out[2]
    PORT
      LAYER met2 ;
        RECT 38.730 0.000 39.010 4.000 ;
    END
  END chany_bottom_out[2]
  PIN chany_bottom_out[3]
    PORT
      LAYER met2 ;
        RECT 29.070 96.000 29.350 100.000 ;
    END
  END chany_bottom_out[3]
  PIN chany_bottom_out[4]
    PORT
      LAYER met3 ;
        RECT 96.000 95.240 100.000 95.840 ;
    END
  END chany_bottom_out[4]
  PIN chany_bottom_out[5]
    PORT
      LAYER met2 ;
        RECT 61.270 96.000 61.550 100.000 ;
    END
  END chany_bottom_out[5]
  PIN chany_bottom_out[6]
    PORT
      LAYER met3 ;
        RECT 0.000 98.640 4.000 99.240 ;
    END
  END chany_bottom_out[6]
  PIN chany_bottom_out[7]
    PORT
      LAYER met2 ;
        RECT 70.930 96.000 71.210 100.000 ;
    END
  END chany_bottom_out[7]
  PIN chany_bottom_out[8]
    PORT
      LAYER met2 ;
        RECT 45.170 96.000 45.450 100.000 ;
    END
  END chany_bottom_out[8]
  PIN chany_bottom_out[9]
    PORT
      LAYER met3 ;
        RECT 96.000 78.240 100.000 78.840 ;
    END
  END chany_bottom_out[9]
  PIN chany_top_in[0]
    PORT
      LAYER met3 ;
        RECT 96.000 61.240 100.000 61.840 ;
    END
  END chany_top_in[0]
  PIN chany_top_in[10]
    PORT
      LAYER met3 ;
        RECT 0.000 6.840 4.000 7.440 ;
    END
  END chany_top_in[10]
  PIN chany_top_in[1]
    PORT
      LAYER met2 ;
        RECT 87.030 96.000 87.310 100.000 ;
    END
  END chany_top_in[1]
  PIN chany_top_in[2]
    PORT
      LAYER met2 ;
        RECT 6.530 0.000 6.810 4.000 ;
    END
  END chany_top_in[2]
  PIN chany_top_in[3]
    PORT
      LAYER met2 ;
        RECT 0.090 0.000 0.370 4.000 ;
    END
  END chany_top_in[3]
  PIN chany_top_in[4]
    PORT
      LAYER met3 ;
        RECT 0.000 23.840 4.000 24.440 ;
    END
  END chany_top_in[4]
  PIN chany_top_in[5]
    PORT
      LAYER met3 ;
        RECT 96.000 71.440 100.000 72.040 ;
    END
  END chany_top_in[5]
  PIN chany_top_in[6]
    PORT
      LAYER met2 ;
        RECT 29.070 0.000 29.350 4.000 ;
    END
  END chany_top_in[6]
  PIN chany_top_in[7]
    PORT
      LAYER met3 ;
        RECT 96.000 54.440 100.000 55.040 ;
    END
  END chany_top_in[7]
  PIN chany_top_in[8]
    PORT
      LAYER met2 ;
        RECT 87.030 0.000 87.310 4.000 ;
    END
  END chany_top_in[8]
  PIN chany_top_in[9]
    PORT
      LAYER met2 ;
        RECT 54.830 96.000 55.110 100.000 ;
    END
  END chany_top_in[9]
  PIN chany_top_out[0]
    PORT
      LAYER met3 ;
        RECT 96.000 27.240 100.000 27.840 ;
    END
  END chany_top_out[0]
  PIN chany_top_out[10]
    PORT
      LAYER met2 ;
        RECT 12.970 0.000 13.250 4.000 ;
    END
  END chany_top_out[10]
  PIN chany_top_out[1]
    PORT
      LAYER met2 ;
        RECT 22.630 0.000 22.910 4.000 ;
    END
  END chany_top_out[1]
  PIN chany_top_out[2]
    PORT
      LAYER met3 ;
        RECT 0.000 74.840 4.000 75.440 ;
    END
  END chany_top_out[2]
  PIN chany_top_out[3]
    PORT
      LAYER met3 ;
        RECT 96.000 37.440 100.000 38.040 ;
    END
  END chany_top_out[3]
  PIN chany_top_out[4]
    PORT
      LAYER met2 ;
        RECT 45.170 0.000 45.450 4.000 ;
    END
  END chany_top_out[4]
  PIN chany_top_out[5]
    PORT
      LAYER met3 ;
        RECT 0.000 57.840 4.000 58.440 ;
    END
  END chany_top_out[5]
  PIN chany_top_out[6]
    PORT
      LAYER met2 ;
        RECT 93.470 96.000 93.750 100.000 ;
    END
  END chany_top_out[6]
  PIN chany_top_out[7]
    PORT
      LAYER met2 ;
        RECT 22.630 96.000 22.910 100.000 ;
    END
  END chany_top_out[7]
  PIN chany_top_out[8]
    PORT
      LAYER met2 ;
        RECT 38.730 96.000 39.010 100.000 ;
    END
  END chany_top_out[8]
  PIN chany_top_out[9]
    PORT
      LAYER met2 ;
        RECT 61.270 0.000 61.550 4.000 ;
    END
  END chany_top_out[9]
  PIN left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_
    PORT
      LAYER met3 ;
        RECT 0.000 40.840 4.000 41.440 ;
    END
  END left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_
  PIN prog_clk
    PORT
      LAYER met3 ;
        RECT 0.000 91.840 4.000 92.440 ;
    END
  END prog_clk
  PIN right_grid_left_width_0_height_0_subtile_0__pin_clk_0_
    PORT
      LAYER met3 ;
        RECT 96.000 44.240 100.000 44.840 ;
    END
  END right_grid_left_width_0_height_0_subtile_0__pin_clk_0_
  PIN vccd1
    PORT
      LAYER met4 ;
        RECT 82.400 10.640 84.000 87.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 60.205 10.640 61.805 87.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 38.010 10.640 39.610 87.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 15.815 10.640 17.415 87.280 ;
    END
  END vccd1
  PIN vssd1
    PORT
      LAYER met4 ;
        RECT 93.495 10.640 95.095 87.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 71.300 10.640 72.900 87.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 49.105 10.640 50.705 87.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 26.910 10.640 28.510 87.280 ;
    END
  END vssd1
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 94.300 87.125 ;
      LAYER met1 ;
        RECT 0.070 10.640 96.070 87.280 ;
      LAYER met2 ;
        RECT 0.100 95.720 6.250 99.125 ;
        RECT 7.090 95.720 12.690 99.125 ;
        RECT 13.530 95.720 22.350 99.125 ;
        RECT 23.190 95.720 28.790 99.125 ;
        RECT 29.630 95.720 38.450 99.125 ;
        RECT 39.290 95.720 44.890 99.125 ;
        RECT 45.730 95.720 54.550 99.125 ;
        RECT 55.390 95.720 60.990 99.125 ;
        RECT 61.830 95.720 70.650 99.125 ;
        RECT 71.490 95.720 77.090 99.125 ;
        RECT 77.930 95.720 86.750 99.125 ;
        RECT 87.590 95.720 93.190 99.125 ;
        RECT 94.030 95.720 96.050 99.125 ;
        RECT 0.100 4.280 96.050 95.720 ;
        RECT 0.650 3.555 6.250 4.280 ;
        RECT 7.090 3.555 12.690 4.280 ;
        RECT 13.530 3.555 22.350 4.280 ;
        RECT 23.190 3.555 28.790 4.280 ;
        RECT 29.630 3.555 38.450 4.280 ;
        RECT 39.290 3.555 44.890 4.280 ;
        RECT 45.730 3.555 54.550 4.280 ;
        RECT 55.390 3.555 60.990 4.280 ;
        RECT 61.830 3.555 70.650 4.280 ;
        RECT 71.490 3.555 77.090 4.280 ;
        RECT 77.930 3.555 86.750 4.280 ;
        RECT 87.590 3.555 93.190 4.280 ;
        RECT 94.030 3.555 96.050 4.280 ;
      LAYER met3 ;
        RECT 4.400 98.240 96.060 99.105 ;
        RECT 4.000 96.240 96.060 98.240 ;
        RECT 4.000 94.840 95.600 96.240 ;
        RECT 4.000 92.840 96.060 94.840 ;
        RECT 4.400 91.440 96.060 92.840 ;
        RECT 4.000 89.440 96.060 91.440 ;
        RECT 4.000 88.040 95.600 89.440 ;
        RECT 4.000 82.640 96.060 88.040 ;
        RECT 4.400 81.240 96.060 82.640 ;
        RECT 4.000 79.240 96.060 81.240 ;
        RECT 4.000 77.840 95.600 79.240 ;
        RECT 4.000 75.840 96.060 77.840 ;
        RECT 4.400 74.440 96.060 75.840 ;
        RECT 4.000 72.440 96.060 74.440 ;
        RECT 4.000 71.040 95.600 72.440 ;
        RECT 4.000 65.640 96.060 71.040 ;
        RECT 4.400 64.240 96.060 65.640 ;
        RECT 4.000 62.240 96.060 64.240 ;
        RECT 4.000 60.840 95.600 62.240 ;
        RECT 4.000 58.840 96.060 60.840 ;
        RECT 4.400 57.440 96.060 58.840 ;
        RECT 4.000 55.440 96.060 57.440 ;
        RECT 4.000 54.040 95.600 55.440 ;
        RECT 4.000 48.640 96.060 54.040 ;
        RECT 4.400 47.240 96.060 48.640 ;
        RECT 4.000 45.240 96.060 47.240 ;
        RECT 4.000 43.840 95.600 45.240 ;
        RECT 4.000 41.840 96.060 43.840 ;
        RECT 4.400 40.440 96.060 41.840 ;
        RECT 4.000 38.440 96.060 40.440 ;
        RECT 4.000 37.040 95.600 38.440 ;
        RECT 4.000 31.640 96.060 37.040 ;
        RECT 4.400 30.240 96.060 31.640 ;
        RECT 4.000 28.240 96.060 30.240 ;
        RECT 4.000 26.840 95.600 28.240 ;
        RECT 4.000 24.840 96.060 26.840 ;
        RECT 4.400 23.440 96.060 24.840 ;
        RECT 4.000 21.440 96.060 23.440 ;
        RECT 4.000 20.040 95.600 21.440 ;
        RECT 4.000 14.640 96.060 20.040 ;
        RECT 4.400 13.240 96.060 14.640 ;
        RECT 4.000 11.240 96.060 13.240 ;
        RECT 4.000 9.840 95.600 11.240 ;
        RECT 4.000 7.840 96.060 9.840 ;
        RECT 4.400 6.440 96.060 7.840 ;
        RECT 4.000 4.440 96.060 6.440 ;
        RECT 4.000 3.575 95.600 4.440 ;
  END
END cby_0__1_
END LIBRARY

