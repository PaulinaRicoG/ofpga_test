VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO user_proj_example
  CLASS BLOCK ;
  FOREIGN user_proj_example ;
  ORIGIN 0.000 0.000 ;
  SIZE 2100.000 BY 3300.000 ;
  PIN io_in[0]
    PORT
      LAYER met3 ;
        RECT 2096.000 69.400 2100.000 70.000 ;
    END
  END io_in[0]
  PIN io_in[10]
    PORT
      LAYER met3 ;
        RECT 0.000 2404.520 4.000 2405.120 ;
    END
  END io_in[10]
  PIN io_in[11]
    PORT
      LAYER met3 ;
        RECT 0.000 1992.440 4.000 1993.040 ;
    END
  END io_in[11]
  PIN io_in[12]
    PORT
      LAYER met3 ;
        RECT 0.000 1580.360 4.000 1580.960 ;
    END
  END io_in[12]
  PIN io_in[13]
    PORT
      LAYER met3 ;
        RECT 0.000 1168.280 4.000 1168.880 ;
    END
  END io_in[13]
  PIN io_in[14]
    PORT
      LAYER met3 ;
        RECT 0.000 756.200 4.000 756.800 ;
    END
  END io_in[14]
  PIN io_in[15]
    PORT
      LAYER met3 ;
        RECT 0.000 344.120 4.000 344.720 ;
    END
  END io_in[15]
  PIN io_in[1]
    PORT
      LAYER met3 ;
        RECT 2096.000 481.480 2100.000 482.080 ;
    END
  END io_in[1]
  PIN io_in[2]
    PORT
      LAYER met3 ;
        RECT 2096.000 893.560 2100.000 894.160 ;
    END
  END io_in[2]
  PIN io_in[3]
    PORT
      LAYER met3 ;
        RECT 2096.000 1305.640 2100.000 1306.240 ;
    END
  END io_in[3]
  PIN io_in[4]
    PORT
      LAYER met3 ;
        RECT 2096.000 1717.720 2100.000 1718.320 ;
    END
  END io_in[4]
  PIN io_in[5]
    PORT
      LAYER met3 ;
        RECT 2096.000 2129.800 2100.000 2130.400 ;
    END
  END io_in[5]
  PIN io_in[6]
    PORT
      LAYER met3 ;
        RECT 2096.000 2541.880 2100.000 2542.480 ;
    END
  END io_in[6]
  PIN io_in[7]
    PORT
      LAYER met3 ;
        RECT 2096.000 2953.960 2100.000 2954.560 ;
    END
  END io_in[7]
  PIN io_in[8]
    PORT
      LAYER met3 ;
        RECT 0.000 3228.680 4.000 3229.280 ;
    END
  END io_in[8]
  PIN io_in[9]
    PORT
      LAYER met3 ;
        RECT 0.000 2816.600 4.000 2817.200 ;
    END
  END io_in[9]
  PIN io_oeb[0]
    PORT
      LAYER met3 ;
        RECT 2096.000 344.120 2100.000 344.720 ;
    END
  END io_oeb[0]
  PIN io_oeb[10]
    PORT
      LAYER met3 ;
        RECT 0.000 2129.800 4.000 2130.400 ;
    END
  END io_oeb[10]
  PIN io_oeb[11]
    PORT
      LAYER met3 ;
        RECT 0.000 1717.720 4.000 1718.320 ;
    END
  END io_oeb[11]
  PIN io_oeb[12]
    PORT
      LAYER met3 ;
        RECT 0.000 1305.640 4.000 1306.240 ;
    END
  END io_oeb[12]
  PIN io_oeb[13]
    PORT
      LAYER met3 ;
        RECT 0.000 893.560 4.000 894.160 ;
    END
  END io_oeb[13]
  PIN io_oeb[14]
    PORT
      LAYER met3 ;
        RECT 0.000 481.480 4.000 482.080 ;
    END
  END io_oeb[14]
  PIN io_oeb[15]
    PORT
      LAYER met3 ;
        RECT 0.000 69.400 4.000 70.000 ;
    END
  END io_oeb[15]
  PIN io_oeb[1]
    PORT
      LAYER met3 ;
        RECT 2096.000 756.200 2100.000 756.800 ;
    END
  END io_oeb[1]
  PIN io_oeb[2]
    PORT
      LAYER met3 ;
        RECT 2096.000 1168.280 2100.000 1168.880 ;
    END
  END io_oeb[2]
  PIN io_oeb[3]
    PORT
      LAYER met3 ;
        RECT 2096.000 1580.360 2100.000 1580.960 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    PORT
      LAYER met3 ;
        RECT 2096.000 1992.440 2100.000 1993.040 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    PORT
      LAYER met3 ;
        RECT 2096.000 2404.520 2100.000 2405.120 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    PORT
      LAYER met3 ;
        RECT 2096.000 2816.600 2100.000 2817.200 ;
    END
  END io_oeb[6]
  PIN io_oeb[7]
    PORT
      LAYER met3 ;
        RECT 2096.000 3228.680 2100.000 3229.280 ;
    END
  END io_oeb[7]
  PIN io_oeb[8]
    PORT
      LAYER met3 ;
        RECT 0.000 2953.960 4.000 2954.560 ;
    END
  END io_oeb[8]
  PIN io_oeb[9]
    PORT
      LAYER met3 ;
        RECT 0.000 2541.880 4.000 2542.480 ;
    END
  END io_oeb[9]
  PIN io_out[0]
    PORT
      LAYER met3 ;
        RECT 2096.000 206.760 2100.000 207.360 ;
    END
  END io_out[0]
  PIN io_out[10]
    PORT
      LAYER met3 ;
        RECT 0.000 2267.160 4.000 2267.760 ;
    END
  END io_out[10]
  PIN io_out[11]
    PORT
      LAYER met3 ;
        RECT 0.000 1855.080 4.000 1855.680 ;
    END
  END io_out[11]
  PIN io_out[12]
    PORT
      LAYER met3 ;
        RECT 0.000 1443.000 4.000 1443.600 ;
    END
  END io_out[12]
  PIN io_out[13]
    PORT
      LAYER met3 ;
        RECT 0.000 1030.920 4.000 1031.520 ;
    END
  END io_out[13]
  PIN io_out[14]
    PORT
      LAYER met3 ;
        RECT 0.000 618.840 4.000 619.440 ;
    END
  END io_out[14]
  PIN io_out[15]
    PORT
      LAYER met3 ;
        RECT 0.000 206.760 4.000 207.360 ;
    END
  END io_out[15]
  PIN io_out[1]
    PORT
      LAYER met3 ;
        RECT 2096.000 618.840 2100.000 619.440 ;
    END
  END io_out[1]
  PIN io_out[2]
    PORT
      LAYER met3 ;
        RECT 2096.000 1030.920 2100.000 1031.520 ;
    END
  END io_out[2]
  PIN io_out[3]
    PORT
      LAYER met3 ;
        RECT 2096.000 1443.000 2100.000 1443.600 ;
    END
  END io_out[3]
  PIN io_out[4]
    PORT
      LAYER met3 ;
        RECT 2096.000 1855.080 2100.000 1855.680 ;
    END
  END io_out[4]
  PIN io_out[5]
    PORT
      LAYER met3 ;
        RECT 2096.000 2267.160 2100.000 2267.760 ;
    END
  END io_out[5]
  PIN io_out[6]
    PORT
      LAYER met3 ;
        RECT 2096.000 2679.240 2100.000 2679.840 ;
    END
  END io_out[6]
  PIN io_out[7]
    PORT
      LAYER met3 ;
        RECT 2096.000 3091.320 2100.000 3091.920 ;
    END
  END io_out[7]
  PIN io_out[8]
    PORT
      LAYER met3 ;
        RECT 0.000 3091.320 4.000 3091.920 ;
    END
  END io_out[8]
  PIN io_out[9]
    PORT
      LAYER met3 ;
        RECT 0.000 2679.240 4.000 2679.840 ;
    END
  END io_out[9]
  PIN irq[0]
    PORT
      LAYER met2 ;
        RECT 2016.270 3296.000 2016.550 3300.000 ;
    END
  END irq[0]
  PIN irq[1]
    PORT
      LAYER met2 ;
        RECT 2021.330 3296.000 2021.610 3300.000 ;
    END
  END irq[1]
  PIN irq[2]
    PORT
      LAYER met2 ;
        RECT 2026.390 3296.000 2026.670 3300.000 ;
    END
  END irq[2]
  PIN la_data_in[0]
    PORT
      LAYER met2 ;
        RECT 73.230 3296.000 73.510 3300.000 ;
    END
  END la_data_in[0]
  PIN la_data_in[100]
    PORT
      LAYER met2 ;
        RECT 1591.230 3296.000 1591.510 3300.000 ;
    END
  END la_data_in[100]
  PIN la_data_in[101]
    PORT
      LAYER met2 ;
        RECT 1606.410 3296.000 1606.690 3300.000 ;
    END
  END la_data_in[101]
  PIN la_data_in[102]
    PORT
      LAYER met2 ;
        RECT 1621.590 3296.000 1621.870 3300.000 ;
    END
  END la_data_in[102]
  PIN la_data_in[103]
    PORT
      LAYER met2 ;
        RECT 1636.770 3296.000 1637.050 3300.000 ;
    END
  END la_data_in[103]
  PIN la_data_in[104]
    PORT
      LAYER met2 ;
        RECT 1651.950 3296.000 1652.230 3300.000 ;
    END
  END la_data_in[104]
  PIN la_data_in[105]
    PORT
      LAYER met2 ;
        RECT 1667.130 3296.000 1667.410 3300.000 ;
    END
  END la_data_in[105]
  PIN la_data_in[106]
    PORT
      LAYER met2 ;
        RECT 1682.310 3296.000 1682.590 3300.000 ;
    END
  END la_data_in[106]
  PIN la_data_in[107]
    PORT
      LAYER met2 ;
        RECT 1697.490 3296.000 1697.770 3300.000 ;
    END
  END la_data_in[107]
  PIN la_data_in[108]
    PORT
      LAYER met2 ;
        RECT 1712.670 3296.000 1712.950 3300.000 ;
    END
  END la_data_in[108]
  PIN la_data_in[109]
    PORT
      LAYER met2 ;
        RECT 1727.850 3296.000 1728.130 3300.000 ;
    END
  END la_data_in[109]
  PIN la_data_in[10]
    PORT
      LAYER met2 ;
        RECT 225.030 3296.000 225.310 3300.000 ;
    END
  END la_data_in[10]
  PIN la_data_in[110]
    PORT
      LAYER met2 ;
        RECT 1743.030 3296.000 1743.310 3300.000 ;
    END
  END la_data_in[110]
  PIN la_data_in[111]
    PORT
      LAYER met2 ;
        RECT 1758.210 3296.000 1758.490 3300.000 ;
    END
  END la_data_in[111]
  PIN la_data_in[112]
    PORT
      LAYER met2 ;
        RECT 1773.390 3296.000 1773.670 3300.000 ;
    END
  END la_data_in[112]
  PIN la_data_in[113]
    PORT
      LAYER met2 ;
        RECT 1788.570 3296.000 1788.850 3300.000 ;
    END
  END la_data_in[113]
  PIN la_data_in[114]
    PORT
      LAYER met2 ;
        RECT 1803.750 3296.000 1804.030 3300.000 ;
    END
  END la_data_in[114]
  PIN la_data_in[115]
    PORT
      LAYER met2 ;
        RECT 1818.930 3296.000 1819.210 3300.000 ;
    END
  END la_data_in[115]
  PIN la_data_in[116]
    PORT
      LAYER met2 ;
        RECT 1834.110 3296.000 1834.390 3300.000 ;
    END
  END la_data_in[116]
  PIN la_data_in[117]
    PORT
      LAYER met2 ;
        RECT 1849.290 3296.000 1849.570 3300.000 ;
    END
  END la_data_in[117]
  PIN la_data_in[118]
    PORT
      LAYER met2 ;
        RECT 1864.470 3296.000 1864.750 3300.000 ;
    END
  END la_data_in[118]
  PIN la_data_in[119]
    PORT
      LAYER met2 ;
        RECT 1879.650 3296.000 1879.930 3300.000 ;
    END
  END la_data_in[119]
  PIN la_data_in[11]
    PORT
      LAYER met2 ;
        RECT 240.210 3296.000 240.490 3300.000 ;
    END
  END la_data_in[11]
  PIN la_data_in[120]
    PORT
      LAYER met2 ;
        RECT 1894.830 3296.000 1895.110 3300.000 ;
    END
  END la_data_in[120]
  PIN la_data_in[121]
    PORT
      LAYER met2 ;
        RECT 1910.010 3296.000 1910.290 3300.000 ;
    END
  END la_data_in[121]
  PIN la_data_in[122]
    PORT
      LAYER met2 ;
        RECT 1925.190 3296.000 1925.470 3300.000 ;
    END
  END la_data_in[122]
  PIN la_data_in[123]
    PORT
      LAYER met2 ;
        RECT 1940.370 3296.000 1940.650 3300.000 ;
    END
  END la_data_in[123]
  PIN la_data_in[124]
    PORT
      LAYER met2 ;
        RECT 1955.550 3296.000 1955.830 3300.000 ;
    END
  END la_data_in[124]
  PIN la_data_in[125]
    PORT
      LAYER met2 ;
        RECT 1970.730 3296.000 1971.010 3300.000 ;
    END
  END la_data_in[125]
  PIN la_data_in[126]
    PORT
      LAYER met2 ;
        RECT 1985.910 3296.000 1986.190 3300.000 ;
    END
  END la_data_in[126]
  PIN la_data_in[127]
    PORT
      LAYER met2 ;
        RECT 2001.090 3296.000 2001.370 3300.000 ;
    END
  END la_data_in[127]
  PIN la_data_in[12]
    PORT
      LAYER met2 ;
        RECT 255.390 3296.000 255.670 3300.000 ;
    END
  END la_data_in[12]
  PIN la_data_in[13]
    PORT
      LAYER met2 ;
        RECT 270.570 3296.000 270.850 3300.000 ;
    END
  END la_data_in[13]
  PIN la_data_in[14]
    PORT
      LAYER met2 ;
        RECT 285.750 3296.000 286.030 3300.000 ;
    END
  END la_data_in[14]
  PIN la_data_in[15]
    PORT
      LAYER met2 ;
        RECT 300.930 3296.000 301.210 3300.000 ;
    END
  END la_data_in[15]
  PIN la_data_in[16]
    PORT
      LAYER met2 ;
        RECT 316.110 3296.000 316.390 3300.000 ;
    END
  END la_data_in[16]
  PIN la_data_in[17]
    PORT
      LAYER met2 ;
        RECT 331.290 3296.000 331.570 3300.000 ;
    END
  END la_data_in[17]
  PIN la_data_in[18]
    PORT
      LAYER met2 ;
        RECT 346.470 3296.000 346.750 3300.000 ;
    END
  END la_data_in[18]
  PIN la_data_in[19]
    PORT
      LAYER met2 ;
        RECT 361.650 3296.000 361.930 3300.000 ;
    END
  END la_data_in[19]
  PIN la_data_in[1]
    PORT
      LAYER met2 ;
        RECT 88.410 3296.000 88.690 3300.000 ;
    END
  END la_data_in[1]
  PIN la_data_in[20]
    PORT
      LAYER met2 ;
        RECT 376.830 3296.000 377.110 3300.000 ;
    END
  END la_data_in[20]
  PIN la_data_in[21]
    PORT
      LAYER met2 ;
        RECT 392.010 3296.000 392.290 3300.000 ;
    END
  END la_data_in[21]
  PIN la_data_in[22]
    PORT
      LAYER met2 ;
        RECT 407.190 3296.000 407.470 3300.000 ;
    END
  END la_data_in[22]
  PIN la_data_in[23]
    PORT
      LAYER met2 ;
        RECT 422.370 3296.000 422.650 3300.000 ;
    END
  END la_data_in[23]
  PIN la_data_in[24]
    PORT
      LAYER met2 ;
        RECT 437.550 3296.000 437.830 3300.000 ;
    END
  END la_data_in[24]
  PIN la_data_in[25]
    PORT
      LAYER met2 ;
        RECT 452.730 3296.000 453.010 3300.000 ;
    END
  END la_data_in[25]
  PIN la_data_in[26]
    PORT
      LAYER met2 ;
        RECT 467.910 3296.000 468.190 3300.000 ;
    END
  END la_data_in[26]
  PIN la_data_in[27]
    PORT
      LAYER met2 ;
        RECT 483.090 3296.000 483.370 3300.000 ;
    END
  END la_data_in[27]
  PIN la_data_in[28]
    PORT
      LAYER met2 ;
        RECT 498.270 3296.000 498.550 3300.000 ;
    END
  END la_data_in[28]
  PIN la_data_in[29]
    PORT
      LAYER met2 ;
        RECT 513.450 3296.000 513.730 3300.000 ;
    END
  END la_data_in[29]
  PIN la_data_in[2]
    PORT
      LAYER met2 ;
        RECT 103.590 3296.000 103.870 3300.000 ;
    END
  END la_data_in[2]
  PIN la_data_in[30]
    PORT
      LAYER met2 ;
        RECT 528.630 3296.000 528.910 3300.000 ;
    END
  END la_data_in[30]
  PIN la_data_in[31]
    PORT
      LAYER met2 ;
        RECT 543.810 3296.000 544.090 3300.000 ;
    END
  END la_data_in[31]
  PIN la_data_in[32]
    PORT
      LAYER met2 ;
        RECT 558.990 3296.000 559.270 3300.000 ;
    END
  END la_data_in[32]
  PIN la_data_in[33]
    PORT
      LAYER met2 ;
        RECT 574.170 3296.000 574.450 3300.000 ;
    END
  END la_data_in[33]
  PIN la_data_in[34]
    PORT
      LAYER met2 ;
        RECT 589.350 3296.000 589.630 3300.000 ;
    END
  END la_data_in[34]
  PIN la_data_in[35]
    PORT
      LAYER met2 ;
        RECT 604.530 3296.000 604.810 3300.000 ;
    END
  END la_data_in[35]
  PIN la_data_in[36]
    PORT
      LAYER met2 ;
        RECT 619.710 3296.000 619.990 3300.000 ;
    END
  END la_data_in[36]
  PIN la_data_in[37]
    PORT
      LAYER met2 ;
        RECT 634.890 3296.000 635.170 3300.000 ;
    END
  END la_data_in[37]
  PIN la_data_in[38]
    PORT
      LAYER met2 ;
        RECT 650.070 3296.000 650.350 3300.000 ;
    END
  END la_data_in[38]
  PIN la_data_in[39]
    PORT
      LAYER met2 ;
        RECT 665.250 3296.000 665.530 3300.000 ;
    END
  END la_data_in[39]
  PIN la_data_in[3]
    PORT
      LAYER met2 ;
        RECT 118.770 3296.000 119.050 3300.000 ;
    END
  END la_data_in[3]
  PIN la_data_in[40]
    PORT
      LAYER met2 ;
        RECT 680.430 3296.000 680.710 3300.000 ;
    END
  END la_data_in[40]
  PIN la_data_in[41]
    PORT
      LAYER met2 ;
        RECT 695.610 3296.000 695.890 3300.000 ;
    END
  END la_data_in[41]
  PIN la_data_in[42]
    PORT
      LAYER met2 ;
        RECT 710.790 3296.000 711.070 3300.000 ;
    END
  END la_data_in[42]
  PIN la_data_in[43]
    PORT
      LAYER met2 ;
        RECT 725.970 3296.000 726.250 3300.000 ;
    END
  END la_data_in[43]
  PIN la_data_in[44]
    PORT
      LAYER met2 ;
        RECT 741.150 3296.000 741.430 3300.000 ;
    END
  END la_data_in[44]
  PIN la_data_in[45]
    PORT
      LAYER met2 ;
        RECT 756.330 3296.000 756.610 3300.000 ;
    END
  END la_data_in[45]
  PIN la_data_in[46]
    PORT
      LAYER met2 ;
        RECT 771.510 3296.000 771.790 3300.000 ;
    END
  END la_data_in[46]
  PIN la_data_in[47]
    PORT
      LAYER met2 ;
        RECT 786.690 3296.000 786.970 3300.000 ;
    END
  END la_data_in[47]
  PIN la_data_in[48]
    PORT
      LAYER met2 ;
        RECT 801.870 3296.000 802.150 3300.000 ;
    END
  END la_data_in[48]
  PIN la_data_in[49]
    PORT
      LAYER met2 ;
        RECT 817.050 3296.000 817.330 3300.000 ;
    END
  END la_data_in[49]
  PIN la_data_in[4]
    PORT
      LAYER met2 ;
        RECT 133.950 3296.000 134.230 3300.000 ;
    END
  END la_data_in[4]
  PIN la_data_in[50]
    PORT
      LAYER met2 ;
        RECT 832.230 3296.000 832.510 3300.000 ;
    END
  END la_data_in[50]
  PIN la_data_in[51]
    PORT
      LAYER met2 ;
        RECT 847.410 3296.000 847.690 3300.000 ;
    END
  END la_data_in[51]
  PIN la_data_in[52]
    PORT
      LAYER met2 ;
        RECT 862.590 3296.000 862.870 3300.000 ;
    END
  END la_data_in[52]
  PIN la_data_in[53]
    PORT
      LAYER met2 ;
        RECT 877.770 3296.000 878.050 3300.000 ;
    END
  END la_data_in[53]
  PIN la_data_in[54]
    PORT
      LAYER met2 ;
        RECT 892.950 3296.000 893.230 3300.000 ;
    END
  END la_data_in[54]
  PIN la_data_in[55]
    PORT
      LAYER met2 ;
        RECT 908.130 3296.000 908.410 3300.000 ;
    END
  END la_data_in[55]
  PIN la_data_in[56]
    PORT
      LAYER met2 ;
        RECT 923.310 3296.000 923.590 3300.000 ;
    END
  END la_data_in[56]
  PIN la_data_in[57]
    PORT
      LAYER met2 ;
        RECT 938.490 3296.000 938.770 3300.000 ;
    END
  END la_data_in[57]
  PIN la_data_in[58]
    PORT
      LAYER met2 ;
        RECT 953.670 3296.000 953.950 3300.000 ;
    END
  END la_data_in[58]
  PIN la_data_in[59]
    PORT
      LAYER met2 ;
        RECT 968.850 3296.000 969.130 3300.000 ;
    END
  END la_data_in[59]
  PIN la_data_in[5]
    PORT
      LAYER met2 ;
        RECT 149.130 3296.000 149.410 3300.000 ;
    END
  END la_data_in[5]
  PIN la_data_in[60]
    PORT
      LAYER met2 ;
        RECT 984.030 3296.000 984.310 3300.000 ;
    END
  END la_data_in[60]
  PIN la_data_in[61]
    PORT
      LAYER met2 ;
        RECT 999.210 3296.000 999.490 3300.000 ;
    END
  END la_data_in[61]
  PIN la_data_in[62]
    PORT
      LAYER met2 ;
        RECT 1014.390 3296.000 1014.670 3300.000 ;
    END
  END la_data_in[62]
  PIN la_data_in[63]
    PORT
      LAYER met2 ;
        RECT 1029.570 3296.000 1029.850 3300.000 ;
    END
  END la_data_in[63]
  PIN la_data_in[64]
    PORT
      LAYER met2 ;
        RECT 1044.750 3296.000 1045.030 3300.000 ;
    END
  END la_data_in[64]
  PIN la_data_in[65]
    PORT
      LAYER met2 ;
        RECT 1059.930 3296.000 1060.210 3300.000 ;
    END
  END la_data_in[65]
  PIN la_data_in[66]
    PORT
      LAYER met2 ;
        RECT 1075.110 3296.000 1075.390 3300.000 ;
    END
  END la_data_in[66]
  PIN la_data_in[67]
    PORT
      LAYER met2 ;
        RECT 1090.290 3296.000 1090.570 3300.000 ;
    END
  END la_data_in[67]
  PIN la_data_in[68]
    PORT
      LAYER met2 ;
        RECT 1105.470 3296.000 1105.750 3300.000 ;
    END
  END la_data_in[68]
  PIN la_data_in[69]
    PORT
      LAYER met2 ;
        RECT 1120.650 3296.000 1120.930 3300.000 ;
    END
  END la_data_in[69]
  PIN la_data_in[6]
    PORT
      LAYER met2 ;
        RECT 164.310 3296.000 164.590 3300.000 ;
    END
  END la_data_in[6]
  PIN la_data_in[70]
    PORT
      LAYER met2 ;
        RECT 1135.830 3296.000 1136.110 3300.000 ;
    END
  END la_data_in[70]
  PIN la_data_in[71]
    PORT
      LAYER met2 ;
        RECT 1151.010 3296.000 1151.290 3300.000 ;
    END
  END la_data_in[71]
  PIN la_data_in[72]
    PORT
      LAYER met2 ;
        RECT 1166.190 3296.000 1166.470 3300.000 ;
    END
  END la_data_in[72]
  PIN la_data_in[73]
    PORT
      LAYER met2 ;
        RECT 1181.370 3296.000 1181.650 3300.000 ;
    END
  END la_data_in[73]
  PIN la_data_in[74]
    PORT
      LAYER met2 ;
        RECT 1196.550 3296.000 1196.830 3300.000 ;
    END
  END la_data_in[74]
  PIN la_data_in[75]
    PORT
      LAYER met2 ;
        RECT 1211.730 3296.000 1212.010 3300.000 ;
    END
  END la_data_in[75]
  PIN la_data_in[76]
    PORT
      LAYER met2 ;
        RECT 1226.910 3296.000 1227.190 3300.000 ;
    END
  END la_data_in[76]
  PIN la_data_in[77]
    PORT
      LAYER met2 ;
        RECT 1242.090 3296.000 1242.370 3300.000 ;
    END
  END la_data_in[77]
  PIN la_data_in[78]
    PORT
      LAYER met2 ;
        RECT 1257.270 3296.000 1257.550 3300.000 ;
    END
  END la_data_in[78]
  PIN la_data_in[79]
    PORT
      LAYER met2 ;
        RECT 1272.450 3296.000 1272.730 3300.000 ;
    END
  END la_data_in[79]
  PIN la_data_in[7]
    PORT
      LAYER met2 ;
        RECT 179.490 3296.000 179.770 3300.000 ;
    END
  END la_data_in[7]
  PIN la_data_in[80]
    PORT
      LAYER met2 ;
        RECT 1287.630 3296.000 1287.910 3300.000 ;
    END
  END la_data_in[80]
  PIN la_data_in[81]
    PORT
      LAYER met2 ;
        RECT 1302.810 3296.000 1303.090 3300.000 ;
    END
  END la_data_in[81]
  PIN la_data_in[82]
    PORT
      LAYER met2 ;
        RECT 1317.990 3296.000 1318.270 3300.000 ;
    END
  END la_data_in[82]
  PIN la_data_in[83]
    PORT
      LAYER met2 ;
        RECT 1333.170 3296.000 1333.450 3300.000 ;
    END
  END la_data_in[83]
  PIN la_data_in[84]
    PORT
      LAYER met2 ;
        RECT 1348.350 3296.000 1348.630 3300.000 ;
    END
  END la_data_in[84]
  PIN la_data_in[85]
    PORT
      LAYER met2 ;
        RECT 1363.530 3296.000 1363.810 3300.000 ;
    END
  END la_data_in[85]
  PIN la_data_in[86]
    PORT
      LAYER met2 ;
        RECT 1378.710 3296.000 1378.990 3300.000 ;
    END
  END la_data_in[86]
  PIN la_data_in[87]
    PORT
      LAYER met2 ;
        RECT 1393.890 3296.000 1394.170 3300.000 ;
    END
  END la_data_in[87]
  PIN la_data_in[88]
    PORT
      LAYER met2 ;
        RECT 1409.070 3296.000 1409.350 3300.000 ;
    END
  END la_data_in[88]
  PIN la_data_in[89]
    PORT
      LAYER met2 ;
        RECT 1424.250 3296.000 1424.530 3300.000 ;
    END
  END la_data_in[89]
  PIN la_data_in[8]
    PORT
      LAYER met2 ;
        RECT 194.670 3296.000 194.950 3300.000 ;
    END
  END la_data_in[8]
  PIN la_data_in[90]
    PORT
      LAYER met2 ;
        RECT 1439.430 3296.000 1439.710 3300.000 ;
    END
  END la_data_in[90]
  PIN la_data_in[91]
    PORT
      LAYER met2 ;
        RECT 1454.610 3296.000 1454.890 3300.000 ;
    END
  END la_data_in[91]
  PIN la_data_in[92]
    PORT
      LAYER met2 ;
        RECT 1469.790 3296.000 1470.070 3300.000 ;
    END
  END la_data_in[92]
  PIN la_data_in[93]
    PORT
      LAYER met2 ;
        RECT 1484.970 3296.000 1485.250 3300.000 ;
    END
  END la_data_in[93]
  PIN la_data_in[94]
    PORT
      LAYER met2 ;
        RECT 1500.150 3296.000 1500.430 3300.000 ;
    END
  END la_data_in[94]
  PIN la_data_in[95]
    PORT
      LAYER met2 ;
        RECT 1515.330 3296.000 1515.610 3300.000 ;
    END
  END la_data_in[95]
  PIN la_data_in[96]
    PORT
      LAYER met2 ;
        RECT 1530.510 3296.000 1530.790 3300.000 ;
    END
  END la_data_in[96]
  PIN la_data_in[97]
    PORT
      LAYER met2 ;
        RECT 1545.690 3296.000 1545.970 3300.000 ;
    END
  END la_data_in[97]
  PIN la_data_in[98]
    PORT
      LAYER met2 ;
        RECT 1560.870 3296.000 1561.150 3300.000 ;
    END
  END la_data_in[98]
  PIN la_data_in[99]
    PORT
      LAYER met2 ;
        RECT 1576.050 3296.000 1576.330 3300.000 ;
    END
  END la_data_in[99]
  PIN la_data_in[9]
    PORT
      LAYER met2 ;
        RECT 209.850 3296.000 210.130 3300.000 ;
    END
  END la_data_in[9]
  PIN la_data_out[0]
    PORT
      LAYER met2 ;
        RECT 78.290 3296.000 78.570 3300.000 ;
    END
  END la_data_out[0]
  PIN la_data_out[100]
    PORT
      LAYER met2 ;
        RECT 1596.290 3296.000 1596.570 3300.000 ;
    END
  END la_data_out[100]
  PIN la_data_out[101]
    PORT
      LAYER met2 ;
        RECT 1611.470 3296.000 1611.750 3300.000 ;
    END
  END la_data_out[101]
  PIN la_data_out[102]
    PORT
      LAYER met2 ;
        RECT 1626.650 3296.000 1626.930 3300.000 ;
    END
  END la_data_out[102]
  PIN la_data_out[103]
    PORT
      LAYER met2 ;
        RECT 1641.830 3296.000 1642.110 3300.000 ;
    END
  END la_data_out[103]
  PIN la_data_out[104]
    PORT
      LAYER met2 ;
        RECT 1657.010 3296.000 1657.290 3300.000 ;
    END
  END la_data_out[104]
  PIN la_data_out[105]
    PORT
      LAYER met2 ;
        RECT 1672.190 3296.000 1672.470 3300.000 ;
    END
  END la_data_out[105]
  PIN la_data_out[106]
    PORT
      LAYER met2 ;
        RECT 1687.370 3296.000 1687.650 3300.000 ;
    END
  END la_data_out[106]
  PIN la_data_out[107]
    PORT
      LAYER met2 ;
        RECT 1702.550 3296.000 1702.830 3300.000 ;
    END
  END la_data_out[107]
  PIN la_data_out[108]
    PORT
      LAYER met2 ;
        RECT 1717.730 3296.000 1718.010 3300.000 ;
    END
  END la_data_out[108]
  PIN la_data_out[109]
    PORT
      LAYER met2 ;
        RECT 1732.910 3296.000 1733.190 3300.000 ;
    END
  END la_data_out[109]
  PIN la_data_out[10]
    PORT
      LAYER met2 ;
        RECT 230.090 3296.000 230.370 3300.000 ;
    END
  END la_data_out[10]
  PIN la_data_out[110]
    PORT
      LAYER met2 ;
        RECT 1748.090 3296.000 1748.370 3300.000 ;
    END
  END la_data_out[110]
  PIN la_data_out[111]
    PORT
      LAYER met2 ;
        RECT 1763.270 3296.000 1763.550 3300.000 ;
    END
  END la_data_out[111]
  PIN la_data_out[112]
    PORT
      LAYER met2 ;
        RECT 1778.450 3296.000 1778.730 3300.000 ;
    END
  END la_data_out[112]
  PIN la_data_out[113]
    PORT
      LAYER met2 ;
        RECT 1793.630 3296.000 1793.910 3300.000 ;
    END
  END la_data_out[113]
  PIN la_data_out[114]
    PORT
      LAYER met2 ;
        RECT 1808.810 3296.000 1809.090 3300.000 ;
    END
  END la_data_out[114]
  PIN la_data_out[115]
    PORT
      LAYER met2 ;
        RECT 1823.990 3296.000 1824.270 3300.000 ;
    END
  END la_data_out[115]
  PIN la_data_out[116]
    PORT
      LAYER met2 ;
        RECT 1839.170 3296.000 1839.450 3300.000 ;
    END
  END la_data_out[116]
  PIN la_data_out[117]
    PORT
      LAYER met2 ;
        RECT 1854.350 3296.000 1854.630 3300.000 ;
    END
  END la_data_out[117]
  PIN la_data_out[118]
    PORT
      LAYER met2 ;
        RECT 1869.530 3296.000 1869.810 3300.000 ;
    END
  END la_data_out[118]
  PIN la_data_out[119]
    PORT
      LAYER met2 ;
        RECT 1884.710 3296.000 1884.990 3300.000 ;
    END
  END la_data_out[119]
  PIN la_data_out[11]
    PORT
      LAYER met2 ;
        RECT 245.270 3296.000 245.550 3300.000 ;
    END
  END la_data_out[11]
  PIN la_data_out[120]
    PORT
      LAYER met2 ;
        RECT 1899.890 3296.000 1900.170 3300.000 ;
    END
  END la_data_out[120]
  PIN la_data_out[121]
    PORT
      LAYER met2 ;
        RECT 1915.070 3296.000 1915.350 3300.000 ;
    END
  END la_data_out[121]
  PIN la_data_out[122]
    PORT
      LAYER met2 ;
        RECT 1930.250 3296.000 1930.530 3300.000 ;
    END
  END la_data_out[122]
  PIN la_data_out[123]
    PORT
      LAYER met2 ;
        RECT 1945.430 3296.000 1945.710 3300.000 ;
    END
  END la_data_out[123]
  PIN la_data_out[124]
    PORT
      LAYER met2 ;
        RECT 1960.610 3296.000 1960.890 3300.000 ;
    END
  END la_data_out[124]
  PIN la_data_out[125]
    PORT
      LAYER met2 ;
        RECT 1975.790 3296.000 1976.070 3300.000 ;
    END
  END la_data_out[125]
  PIN la_data_out[126]
    PORT
      LAYER met2 ;
        RECT 1990.970 3296.000 1991.250 3300.000 ;
    END
  END la_data_out[126]
  PIN la_data_out[127]
    PORT
      LAYER met2 ;
        RECT 2006.150 3296.000 2006.430 3300.000 ;
    END
  END la_data_out[127]
  PIN la_data_out[12]
    PORT
      LAYER met2 ;
        RECT 260.450 3296.000 260.730 3300.000 ;
    END
  END la_data_out[12]
  PIN la_data_out[13]
    PORT
      LAYER met2 ;
        RECT 275.630 3296.000 275.910 3300.000 ;
    END
  END la_data_out[13]
  PIN la_data_out[14]
    PORT
      LAYER met2 ;
        RECT 290.810 3296.000 291.090 3300.000 ;
    END
  END la_data_out[14]
  PIN la_data_out[15]
    PORT
      LAYER met2 ;
        RECT 305.990 3296.000 306.270 3300.000 ;
    END
  END la_data_out[15]
  PIN la_data_out[16]
    PORT
      LAYER met2 ;
        RECT 321.170 3296.000 321.450 3300.000 ;
    END
  END la_data_out[16]
  PIN la_data_out[17]
    PORT
      LAYER met2 ;
        RECT 336.350 3296.000 336.630 3300.000 ;
    END
  END la_data_out[17]
  PIN la_data_out[18]
    PORT
      LAYER met2 ;
        RECT 351.530 3296.000 351.810 3300.000 ;
    END
  END la_data_out[18]
  PIN la_data_out[19]
    PORT
      LAYER met2 ;
        RECT 366.710 3296.000 366.990 3300.000 ;
    END
  END la_data_out[19]
  PIN la_data_out[1]
    PORT
      LAYER met2 ;
        RECT 93.470 3296.000 93.750 3300.000 ;
    END
  END la_data_out[1]
  PIN la_data_out[20]
    PORT
      LAYER met2 ;
        RECT 381.890 3296.000 382.170 3300.000 ;
    END
  END la_data_out[20]
  PIN la_data_out[21]
    PORT
      LAYER met2 ;
        RECT 397.070 3296.000 397.350 3300.000 ;
    END
  END la_data_out[21]
  PIN la_data_out[22]
    PORT
      LAYER met2 ;
        RECT 412.250 3296.000 412.530 3300.000 ;
    END
  END la_data_out[22]
  PIN la_data_out[23]
    PORT
      LAYER met2 ;
        RECT 427.430 3296.000 427.710 3300.000 ;
    END
  END la_data_out[23]
  PIN la_data_out[24]
    PORT
      LAYER met2 ;
        RECT 442.610 3296.000 442.890 3300.000 ;
    END
  END la_data_out[24]
  PIN la_data_out[25]
    PORT
      LAYER met2 ;
        RECT 457.790 3296.000 458.070 3300.000 ;
    END
  END la_data_out[25]
  PIN la_data_out[26]
    PORT
      LAYER met2 ;
        RECT 472.970 3296.000 473.250 3300.000 ;
    END
  END la_data_out[26]
  PIN la_data_out[27]
    PORT
      LAYER met2 ;
        RECT 488.150 3296.000 488.430 3300.000 ;
    END
  END la_data_out[27]
  PIN la_data_out[28]
    PORT
      LAYER met2 ;
        RECT 503.330 3296.000 503.610 3300.000 ;
    END
  END la_data_out[28]
  PIN la_data_out[29]
    PORT
      LAYER met2 ;
        RECT 518.510 3296.000 518.790 3300.000 ;
    END
  END la_data_out[29]
  PIN la_data_out[2]
    PORT
      LAYER met2 ;
        RECT 108.650 3296.000 108.930 3300.000 ;
    END
  END la_data_out[2]
  PIN la_data_out[30]
    PORT
      LAYER met2 ;
        RECT 533.690 3296.000 533.970 3300.000 ;
    END
  END la_data_out[30]
  PIN la_data_out[31]
    PORT
      LAYER met2 ;
        RECT 548.870 3296.000 549.150 3300.000 ;
    END
  END la_data_out[31]
  PIN la_data_out[32]
    PORT
      LAYER met2 ;
        RECT 564.050 3296.000 564.330 3300.000 ;
    END
  END la_data_out[32]
  PIN la_data_out[33]
    PORT
      LAYER met2 ;
        RECT 579.230 3296.000 579.510 3300.000 ;
    END
  END la_data_out[33]
  PIN la_data_out[34]
    PORT
      LAYER met2 ;
        RECT 594.410 3296.000 594.690 3300.000 ;
    END
  END la_data_out[34]
  PIN la_data_out[35]
    PORT
      LAYER met2 ;
        RECT 609.590 3296.000 609.870 3300.000 ;
    END
  END la_data_out[35]
  PIN la_data_out[36]
    PORT
      LAYER met2 ;
        RECT 624.770 3296.000 625.050 3300.000 ;
    END
  END la_data_out[36]
  PIN la_data_out[37]
    PORT
      LAYER met2 ;
        RECT 639.950 3296.000 640.230 3300.000 ;
    END
  END la_data_out[37]
  PIN la_data_out[38]
    PORT
      LAYER met2 ;
        RECT 655.130 3296.000 655.410 3300.000 ;
    END
  END la_data_out[38]
  PIN la_data_out[39]
    PORT
      LAYER met2 ;
        RECT 670.310 3296.000 670.590 3300.000 ;
    END
  END la_data_out[39]
  PIN la_data_out[3]
    PORT
      LAYER met2 ;
        RECT 123.830 3296.000 124.110 3300.000 ;
    END
  END la_data_out[3]
  PIN la_data_out[40]
    PORT
      LAYER met2 ;
        RECT 685.490 3296.000 685.770 3300.000 ;
    END
  END la_data_out[40]
  PIN la_data_out[41]
    PORT
      LAYER met2 ;
        RECT 700.670 3296.000 700.950 3300.000 ;
    END
  END la_data_out[41]
  PIN la_data_out[42]
    PORT
      LAYER met2 ;
        RECT 715.850 3296.000 716.130 3300.000 ;
    END
  END la_data_out[42]
  PIN la_data_out[43]
    PORT
      LAYER met2 ;
        RECT 731.030 3296.000 731.310 3300.000 ;
    END
  END la_data_out[43]
  PIN la_data_out[44]
    PORT
      LAYER met2 ;
        RECT 746.210 3296.000 746.490 3300.000 ;
    END
  END la_data_out[44]
  PIN la_data_out[45]
    PORT
      LAYER met2 ;
        RECT 761.390 3296.000 761.670 3300.000 ;
    END
  END la_data_out[45]
  PIN la_data_out[46]
    PORT
      LAYER met2 ;
        RECT 776.570 3296.000 776.850 3300.000 ;
    END
  END la_data_out[46]
  PIN la_data_out[47]
    PORT
      LAYER met2 ;
        RECT 791.750 3296.000 792.030 3300.000 ;
    END
  END la_data_out[47]
  PIN la_data_out[48]
    PORT
      LAYER met2 ;
        RECT 806.930 3296.000 807.210 3300.000 ;
    END
  END la_data_out[48]
  PIN la_data_out[49]
    PORT
      LAYER met2 ;
        RECT 822.110 3296.000 822.390 3300.000 ;
    END
  END la_data_out[49]
  PIN la_data_out[4]
    PORT
      LAYER met2 ;
        RECT 139.010 3296.000 139.290 3300.000 ;
    END
  END la_data_out[4]
  PIN la_data_out[50]
    PORT
      LAYER met2 ;
        RECT 837.290 3296.000 837.570 3300.000 ;
    END
  END la_data_out[50]
  PIN la_data_out[51]
    PORT
      LAYER met2 ;
        RECT 852.470 3296.000 852.750 3300.000 ;
    END
  END la_data_out[51]
  PIN la_data_out[52]
    PORT
      LAYER met2 ;
        RECT 867.650 3296.000 867.930 3300.000 ;
    END
  END la_data_out[52]
  PIN la_data_out[53]
    PORT
      LAYER met2 ;
        RECT 882.830 3296.000 883.110 3300.000 ;
    END
  END la_data_out[53]
  PIN la_data_out[54]
    PORT
      LAYER met2 ;
        RECT 898.010 3296.000 898.290 3300.000 ;
    END
  END la_data_out[54]
  PIN la_data_out[55]
    PORT
      LAYER met2 ;
        RECT 913.190 3296.000 913.470 3300.000 ;
    END
  END la_data_out[55]
  PIN la_data_out[56]
    PORT
      LAYER met2 ;
        RECT 928.370 3296.000 928.650 3300.000 ;
    END
  END la_data_out[56]
  PIN la_data_out[57]
    PORT
      LAYER met2 ;
        RECT 943.550 3296.000 943.830 3300.000 ;
    END
  END la_data_out[57]
  PIN la_data_out[58]
    PORT
      LAYER met2 ;
        RECT 958.730 3296.000 959.010 3300.000 ;
    END
  END la_data_out[58]
  PIN la_data_out[59]
    PORT
      LAYER met2 ;
        RECT 973.910 3296.000 974.190 3300.000 ;
    END
  END la_data_out[59]
  PIN la_data_out[5]
    PORT
      LAYER met2 ;
        RECT 154.190 3296.000 154.470 3300.000 ;
    END
  END la_data_out[5]
  PIN la_data_out[60]
    PORT
      LAYER met2 ;
        RECT 989.090 3296.000 989.370 3300.000 ;
    END
  END la_data_out[60]
  PIN la_data_out[61]
    PORT
      LAYER met2 ;
        RECT 1004.270 3296.000 1004.550 3300.000 ;
    END
  END la_data_out[61]
  PIN la_data_out[62]
    PORT
      LAYER met2 ;
        RECT 1019.450 3296.000 1019.730 3300.000 ;
    END
  END la_data_out[62]
  PIN la_data_out[63]
    PORT
      LAYER met2 ;
        RECT 1034.630 3296.000 1034.910 3300.000 ;
    END
  END la_data_out[63]
  PIN la_data_out[64]
    PORT
      LAYER met2 ;
        RECT 1049.810 3296.000 1050.090 3300.000 ;
    END
  END la_data_out[64]
  PIN la_data_out[65]
    PORT
      LAYER met2 ;
        RECT 1064.990 3296.000 1065.270 3300.000 ;
    END
  END la_data_out[65]
  PIN la_data_out[66]
    PORT
      LAYER met2 ;
        RECT 1080.170 3296.000 1080.450 3300.000 ;
    END
  END la_data_out[66]
  PIN la_data_out[67]
    PORT
      LAYER met2 ;
        RECT 1095.350 3296.000 1095.630 3300.000 ;
    END
  END la_data_out[67]
  PIN la_data_out[68]
    PORT
      LAYER met2 ;
        RECT 1110.530 3296.000 1110.810 3300.000 ;
    END
  END la_data_out[68]
  PIN la_data_out[69]
    PORT
      LAYER met2 ;
        RECT 1125.710 3296.000 1125.990 3300.000 ;
    END
  END la_data_out[69]
  PIN la_data_out[6]
    PORT
      LAYER met2 ;
        RECT 169.370 3296.000 169.650 3300.000 ;
    END
  END la_data_out[6]
  PIN la_data_out[70]
    PORT
      LAYER met2 ;
        RECT 1140.890 3296.000 1141.170 3300.000 ;
    END
  END la_data_out[70]
  PIN la_data_out[71]
    PORT
      LAYER met2 ;
        RECT 1156.070 3296.000 1156.350 3300.000 ;
    END
  END la_data_out[71]
  PIN la_data_out[72]
    PORT
      LAYER met2 ;
        RECT 1171.250 3296.000 1171.530 3300.000 ;
    END
  END la_data_out[72]
  PIN la_data_out[73]
    PORT
      LAYER met2 ;
        RECT 1186.430 3296.000 1186.710 3300.000 ;
    END
  END la_data_out[73]
  PIN la_data_out[74]
    PORT
      LAYER met2 ;
        RECT 1201.610 3296.000 1201.890 3300.000 ;
    END
  END la_data_out[74]
  PIN la_data_out[75]
    PORT
      LAYER met2 ;
        RECT 1216.790 3296.000 1217.070 3300.000 ;
    END
  END la_data_out[75]
  PIN la_data_out[76]
    PORT
      LAYER met2 ;
        RECT 1231.970 3296.000 1232.250 3300.000 ;
    END
  END la_data_out[76]
  PIN la_data_out[77]
    PORT
      LAYER met2 ;
        RECT 1247.150 3296.000 1247.430 3300.000 ;
    END
  END la_data_out[77]
  PIN la_data_out[78]
    PORT
      LAYER met2 ;
        RECT 1262.330 3296.000 1262.610 3300.000 ;
    END
  END la_data_out[78]
  PIN la_data_out[79]
    PORT
      LAYER met2 ;
        RECT 1277.510 3296.000 1277.790 3300.000 ;
    END
  END la_data_out[79]
  PIN la_data_out[7]
    PORT
      LAYER met2 ;
        RECT 184.550 3296.000 184.830 3300.000 ;
    END
  END la_data_out[7]
  PIN la_data_out[80]
    PORT
      LAYER met2 ;
        RECT 1292.690 3296.000 1292.970 3300.000 ;
    END
  END la_data_out[80]
  PIN la_data_out[81]
    PORT
      LAYER met2 ;
        RECT 1307.870 3296.000 1308.150 3300.000 ;
    END
  END la_data_out[81]
  PIN la_data_out[82]
    PORT
      LAYER met2 ;
        RECT 1323.050 3296.000 1323.330 3300.000 ;
    END
  END la_data_out[82]
  PIN la_data_out[83]
    PORT
      LAYER met2 ;
        RECT 1338.230 3296.000 1338.510 3300.000 ;
    END
  END la_data_out[83]
  PIN la_data_out[84]
    PORT
      LAYER met2 ;
        RECT 1353.410 3296.000 1353.690 3300.000 ;
    END
  END la_data_out[84]
  PIN la_data_out[85]
    PORT
      LAYER met2 ;
        RECT 1368.590 3296.000 1368.870 3300.000 ;
    END
  END la_data_out[85]
  PIN la_data_out[86]
    PORT
      LAYER met2 ;
        RECT 1383.770 3296.000 1384.050 3300.000 ;
    END
  END la_data_out[86]
  PIN la_data_out[87]
    PORT
      LAYER met2 ;
        RECT 1398.950 3296.000 1399.230 3300.000 ;
    END
  END la_data_out[87]
  PIN la_data_out[88]
    PORT
      LAYER met2 ;
        RECT 1414.130 3296.000 1414.410 3300.000 ;
    END
  END la_data_out[88]
  PIN la_data_out[89]
    PORT
      LAYER met2 ;
        RECT 1429.310 3296.000 1429.590 3300.000 ;
    END
  END la_data_out[89]
  PIN la_data_out[8]
    PORT
      LAYER met2 ;
        RECT 199.730 3296.000 200.010 3300.000 ;
    END
  END la_data_out[8]
  PIN la_data_out[90]
    PORT
      LAYER met2 ;
        RECT 1444.490 3296.000 1444.770 3300.000 ;
    END
  END la_data_out[90]
  PIN la_data_out[91]
    PORT
      LAYER met2 ;
        RECT 1459.670 3296.000 1459.950 3300.000 ;
    END
  END la_data_out[91]
  PIN la_data_out[92]
    PORT
      LAYER met2 ;
        RECT 1474.850 3296.000 1475.130 3300.000 ;
    END
  END la_data_out[92]
  PIN la_data_out[93]
    PORT
      LAYER met2 ;
        RECT 1490.030 3296.000 1490.310 3300.000 ;
    END
  END la_data_out[93]
  PIN la_data_out[94]
    PORT
      LAYER met2 ;
        RECT 1505.210 3296.000 1505.490 3300.000 ;
    END
  END la_data_out[94]
  PIN la_data_out[95]
    PORT
      LAYER met2 ;
        RECT 1520.390 3296.000 1520.670 3300.000 ;
    END
  END la_data_out[95]
  PIN la_data_out[96]
    PORT
      LAYER met2 ;
        RECT 1535.570 3296.000 1535.850 3300.000 ;
    END
  END la_data_out[96]
  PIN la_data_out[97]
    PORT
      LAYER met2 ;
        RECT 1550.750 3296.000 1551.030 3300.000 ;
    END
  END la_data_out[97]
  PIN la_data_out[98]
    PORT
      LAYER met2 ;
        RECT 1565.930 3296.000 1566.210 3300.000 ;
    END
  END la_data_out[98]
  PIN la_data_out[99]
    PORT
      LAYER met2 ;
        RECT 1581.110 3296.000 1581.390 3300.000 ;
    END
  END la_data_out[99]
  PIN la_data_out[9]
    PORT
      LAYER met2 ;
        RECT 214.910 3296.000 215.190 3300.000 ;
    END
  END la_data_out[9]
  PIN la_oenb[0]
    PORT
      LAYER met2 ;
        RECT 83.350 3296.000 83.630 3300.000 ;
    END
  END la_oenb[0]
  PIN la_oenb[100]
    PORT
      LAYER met2 ;
        RECT 1601.350 3296.000 1601.630 3300.000 ;
    END
  END la_oenb[100]
  PIN la_oenb[101]
    PORT
      LAYER met2 ;
        RECT 1616.530 3296.000 1616.810 3300.000 ;
    END
  END la_oenb[101]
  PIN la_oenb[102]
    PORT
      LAYER met2 ;
        RECT 1631.710 3296.000 1631.990 3300.000 ;
    END
  END la_oenb[102]
  PIN la_oenb[103]
    PORT
      LAYER met2 ;
        RECT 1646.890 3296.000 1647.170 3300.000 ;
    END
  END la_oenb[103]
  PIN la_oenb[104]
    PORT
      LAYER met2 ;
        RECT 1662.070 3296.000 1662.350 3300.000 ;
    END
  END la_oenb[104]
  PIN la_oenb[105]
    PORT
      LAYER met2 ;
        RECT 1677.250 3296.000 1677.530 3300.000 ;
    END
  END la_oenb[105]
  PIN la_oenb[106]
    PORT
      LAYER met2 ;
        RECT 1692.430 3296.000 1692.710 3300.000 ;
    END
  END la_oenb[106]
  PIN la_oenb[107]
    PORT
      LAYER met2 ;
        RECT 1707.610 3296.000 1707.890 3300.000 ;
    END
  END la_oenb[107]
  PIN la_oenb[108]
    PORT
      LAYER met2 ;
        RECT 1722.790 3296.000 1723.070 3300.000 ;
    END
  END la_oenb[108]
  PIN la_oenb[109]
    PORT
      LAYER met2 ;
        RECT 1737.970 3296.000 1738.250 3300.000 ;
    END
  END la_oenb[109]
  PIN la_oenb[10]
    PORT
      LAYER met2 ;
        RECT 235.150 3296.000 235.430 3300.000 ;
    END
  END la_oenb[10]
  PIN la_oenb[110]
    PORT
      LAYER met2 ;
        RECT 1753.150 3296.000 1753.430 3300.000 ;
    END
  END la_oenb[110]
  PIN la_oenb[111]
    PORT
      LAYER met2 ;
        RECT 1768.330 3296.000 1768.610 3300.000 ;
    END
  END la_oenb[111]
  PIN la_oenb[112]
    PORT
      LAYER met2 ;
        RECT 1783.510 3296.000 1783.790 3300.000 ;
    END
  END la_oenb[112]
  PIN la_oenb[113]
    PORT
      LAYER met2 ;
        RECT 1798.690 3296.000 1798.970 3300.000 ;
    END
  END la_oenb[113]
  PIN la_oenb[114]
    PORT
      LAYER met2 ;
        RECT 1813.870 3296.000 1814.150 3300.000 ;
    END
  END la_oenb[114]
  PIN la_oenb[115]
    PORT
      LAYER met2 ;
        RECT 1829.050 3296.000 1829.330 3300.000 ;
    END
  END la_oenb[115]
  PIN la_oenb[116]
    PORT
      LAYER met2 ;
        RECT 1844.230 3296.000 1844.510 3300.000 ;
    END
  END la_oenb[116]
  PIN la_oenb[117]
    PORT
      LAYER met2 ;
        RECT 1859.410 3296.000 1859.690 3300.000 ;
    END
  END la_oenb[117]
  PIN la_oenb[118]
    PORT
      LAYER met2 ;
        RECT 1874.590 3296.000 1874.870 3300.000 ;
    END
  END la_oenb[118]
  PIN la_oenb[119]
    PORT
      LAYER met2 ;
        RECT 1889.770 3296.000 1890.050 3300.000 ;
    END
  END la_oenb[119]
  PIN la_oenb[11]
    PORT
      LAYER met2 ;
        RECT 250.330 3296.000 250.610 3300.000 ;
    END
  END la_oenb[11]
  PIN la_oenb[120]
    PORT
      LAYER met2 ;
        RECT 1904.950 3296.000 1905.230 3300.000 ;
    END
  END la_oenb[120]
  PIN la_oenb[121]
    PORT
      LAYER met2 ;
        RECT 1920.130 3296.000 1920.410 3300.000 ;
    END
  END la_oenb[121]
  PIN la_oenb[122]
    PORT
      LAYER met2 ;
        RECT 1935.310 3296.000 1935.590 3300.000 ;
    END
  END la_oenb[122]
  PIN la_oenb[123]
    PORT
      LAYER met2 ;
        RECT 1950.490 3296.000 1950.770 3300.000 ;
    END
  END la_oenb[123]
  PIN la_oenb[124]
    PORT
      LAYER met2 ;
        RECT 1965.670 3296.000 1965.950 3300.000 ;
    END
  END la_oenb[124]
  PIN la_oenb[125]
    PORT
      LAYER met2 ;
        RECT 1980.850 3296.000 1981.130 3300.000 ;
    END
  END la_oenb[125]
  PIN la_oenb[126]
    PORT
      LAYER met2 ;
        RECT 1996.030 3296.000 1996.310 3300.000 ;
    END
  END la_oenb[126]
  PIN la_oenb[127]
    PORT
      LAYER met2 ;
        RECT 2011.210 3296.000 2011.490 3300.000 ;
    END
  END la_oenb[127]
  PIN la_oenb[12]
    PORT
      LAYER met2 ;
        RECT 265.510 3296.000 265.790 3300.000 ;
    END
  END la_oenb[12]
  PIN la_oenb[13]
    PORT
      LAYER met2 ;
        RECT 280.690 3296.000 280.970 3300.000 ;
    END
  END la_oenb[13]
  PIN la_oenb[14]
    PORT
      LAYER met2 ;
        RECT 295.870 3296.000 296.150 3300.000 ;
    END
  END la_oenb[14]
  PIN la_oenb[15]
    PORT
      LAYER met2 ;
        RECT 311.050 3296.000 311.330 3300.000 ;
    END
  END la_oenb[15]
  PIN la_oenb[16]
    PORT
      LAYER met2 ;
        RECT 326.230 3296.000 326.510 3300.000 ;
    END
  END la_oenb[16]
  PIN la_oenb[17]
    PORT
      LAYER met2 ;
        RECT 341.410 3296.000 341.690 3300.000 ;
    END
  END la_oenb[17]
  PIN la_oenb[18]
    PORT
      LAYER met2 ;
        RECT 356.590 3296.000 356.870 3300.000 ;
    END
  END la_oenb[18]
  PIN la_oenb[19]
    PORT
      LAYER met2 ;
        RECT 371.770 3296.000 372.050 3300.000 ;
    END
  END la_oenb[19]
  PIN la_oenb[1]
    PORT
      LAYER met2 ;
        RECT 98.530 3296.000 98.810 3300.000 ;
    END
  END la_oenb[1]
  PIN la_oenb[20]
    PORT
      LAYER met2 ;
        RECT 386.950 3296.000 387.230 3300.000 ;
    END
  END la_oenb[20]
  PIN la_oenb[21]
    PORT
      LAYER met2 ;
        RECT 402.130 3296.000 402.410 3300.000 ;
    END
  END la_oenb[21]
  PIN la_oenb[22]
    PORT
      LAYER met2 ;
        RECT 417.310 3296.000 417.590 3300.000 ;
    END
  END la_oenb[22]
  PIN la_oenb[23]
    PORT
      LAYER met2 ;
        RECT 432.490 3296.000 432.770 3300.000 ;
    END
  END la_oenb[23]
  PIN la_oenb[24]
    PORT
      LAYER met2 ;
        RECT 447.670 3296.000 447.950 3300.000 ;
    END
  END la_oenb[24]
  PIN la_oenb[25]
    PORT
      LAYER met2 ;
        RECT 462.850 3296.000 463.130 3300.000 ;
    END
  END la_oenb[25]
  PIN la_oenb[26]
    PORT
      LAYER met2 ;
        RECT 478.030 3296.000 478.310 3300.000 ;
    END
  END la_oenb[26]
  PIN la_oenb[27]
    PORT
      LAYER met2 ;
        RECT 493.210 3296.000 493.490 3300.000 ;
    END
  END la_oenb[27]
  PIN la_oenb[28]
    PORT
      LAYER met2 ;
        RECT 508.390 3296.000 508.670 3300.000 ;
    END
  END la_oenb[28]
  PIN la_oenb[29]
    PORT
      LAYER met2 ;
        RECT 523.570 3296.000 523.850 3300.000 ;
    END
  END la_oenb[29]
  PIN la_oenb[2]
    PORT
      LAYER met2 ;
        RECT 113.710 3296.000 113.990 3300.000 ;
    END
  END la_oenb[2]
  PIN la_oenb[30]
    PORT
      LAYER met2 ;
        RECT 538.750 3296.000 539.030 3300.000 ;
    END
  END la_oenb[30]
  PIN la_oenb[31]
    PORT
      LAYER met2 ;
        RECT 553.930 3296.000 554.210 3300.000 ;
    END
  END la_oenb[31]
  PIN la_oenb[32]
    PORT
      LAYER met2 ;
        RECT 569.110 3296.000 569.390 3300.000 ;
    END
  END la_oenb[32]
  PIN la_oenb[33]
    PORT
      LAYER met2 ;
        RECT 584.290 3296.000 584.570 3300.000 ;
    END
  END la_oenb[33]
  PIN la_oenb[34]
    PORT
      LAYER met2 ;
        RECT 599.470 3296.000 599.750 3300.000 ;
    END
  END la_oenb[34]
  PIN la_oenb[35]
    PORT
      LAYER met2 ;
        RECT 614.650 3296.000 614.930 3300.000 ;
    END
  END la_oenb[35]
  PIN la_oenb[36]
    PORT
      LAYER met2 ;
        RECT 629.830 3296.000 630.110 3300.000 ;
    END
  END la_oenb[36]
  PIN la_oenb[37]
    PORT
      LAYER met2 ;
        RECT 645.010 3296.000 645.290 3300.000 ;
    END
  END la_oenb[37]
  PIN la_oenb[38]
    PORT
      LAYER met2 ;
        RECT 660.190 3296.000 660.470 3300.000 ;
    END
  END la_oenb[38]
  PIN la_oenb[39]
    PORT
      LAYER met2 ;
        RECT 675.370 3296.000 675.650 3300.000 ;
    END
  END la_oenb[39]
  PIN la_oenb[3]
    PORT
      LAYER met2 ;
        RECT 128.890 3296.000 129.170 3300.000 ;
    END
  END la_oenb[3]
  PIN la_oenb[40]
    PORT
      LAYER met2 ;
        RECT 690.550 3296.000 690.830 3300.000 ;
    END
  END la_oenb[40]
  PIN la_oenb[41]
    PORT
      LAYER met2 ;
        RECT 705.730 3296.000 706.010 3300.000 ;
    END
  END la_oenb[41]
  PIN la_oenb[42]
    PORT
      LAYER met2 ;
        RECT 720.910 3296.000 721.190 3300.000 ;
    END
  END la_oenb[42]
  PIN la_oenb[43]
    PORT
      LAYER met2 ;
        RECT 736.090 3296.000 736.370 3300.000 ;
    END
  END la_oenb[43]
  PIN la_oenb[44]
    PORT
      LAYER met2 ;
        RECT 751.270 3296.000 751.550 3300.000 ;
    END
  END la_oenb[44]
  PIN la_oenb[45]
    PORT
      LAYER met2 ;
        RECT 766.450 3296.000 766.730 3300.000 ;
    END
  END la_oenb[45]
  PIN la_oenb[46]
    PORT
      LAYER met2 ;
        RECT 781.630 3296.000 781.910 3300.000 ;
    END
  END la_oenb[46]
  PIN la_oenb[47]
    PORT
      LAYER met2 ;
        RECT 796.810 3296.000 797.090 3300.000 ;
    END
  END la_oenb[47]
  PIN la_oenb[48]
    PORT
      LAYER met2 ;
        RECT 811.990 3296.000 812.270 3300.000 ;
    END
  END la_oenb[48]
  PIN la_oenb[49]
    PORT
      LAYER met2 ;
        RECT 827.170 3296.000 827.450 3300.000 ;
    END
  END la_oenb[49]
  PIN la_oenb[4]
    PORT
      LAYER met2 ;
        RECT 144.070 3296.000 144.350 3300.000 ;
    END
  END la_oenb[4]
  PIN la_oenb[50]
    PORT
      LAYER met2 ;
        RECT 842.350 3296.000 842.630 3300.000 ;
    END
  END la_oenb[50]
  PIN la_oenb[51]
    PORT
      LAYER met2 ;
        RECT 857.530 3296.000 857.810 3300.000 ;
    END
  END la_oenb[51]
  PIN la_oenb[52]
    PORT
      LAYER met2 ;
        RECT 872.710 3296.000 872.990 3300.000 ;
    END
  END la_oenb[52]
  PIN la_oenb[53]
    PORT
      LAYER met2 ;
        RECT 887.890 3296.000 888.170 3300.000 ;
    END
  END la_oenb[53]
  PIN la_oenb[54]
    PORT
      LAYER met2 ;
        RECT 903.070 3296.000 903.350 3300.000 ;
    END
  END la_oenb[54]
  PIN la_oenb[55]
    PORT
      LAYER met2 ;
        RECT 918.250 3296.000 918.530 3300.000 ;
    END
  END la_oenb[55]
  PIN la_oenb[56]
    PORT
      LAYER met2 ;
        RECT 933.430 3296.000 933.710 3300.000 ;
    END
  END la_oenb[56]
  PIN la_oenb[57]
    PORT
      LAYER met2 ;
        RECT 948.610 3296.000 948.890 3300.000 ;
    END
  END la_oenb[57]
  PIN la_oenb[58]
    PORT
      LAYER met2 ;
        RECT 963.790 3296.000 964.070 3300.000 ;
    END
  END la_oenb[58]
  PIN la_oenb[59]
    PORT
      LAYER met2 ;
        RECT 978.970 3296.000 979.250 3300.000 ;
    END
  END la_oenb[59]
  PIN la_oenb[5]
    PORT
      LAYER met2 ;
        RECT 159.250 3296.000 159.530 3300.000 ;
    END
  END la_oenb[5]
  PIN la_oenb[60]
    PORT
      LAYER met2 ;
        RECT 994.150 3296.000 994.430 3300.000 ;
    END
  END la_oenb[60]
  PIN la_oenb[61]
    PORT
      LAYER met2 ;
        RECT 1009.330 3296.000 1009.610 3300.000 ;
    END
  END la_oenb[61]
  PIN la_oenb[62]
    PORT
      LAYER met2 ;
        RECT 1024.510 3296.000 1024.790 3300.000 ;
    END
  END la_oenb[62]
  PIN la_oenb[63]
    PORT
      LAYER met2 ;
        RECT 1039.690 3296.000 1039.970 3300.000 ;
    END
  END la_oenb[63]
  PIN la_oenb[64]
    PORT
      LAYER met2 ;
        RECT 1054.870 3296.000 1055.150 3300.000 ;
    END
  END la_oenb[64]
  PIN la_oenb[65]
    PORT
      LAYER met2 ;
        RECT 1070.050 3296.000 1070.330 3300.000 ;
    END
  END la_oenb[65]
  PIN la_oenb[66]
    PORT
      LAYER met2 ;
        RECT 1085.230 3296.000 1085.510 3300.000 ;
    END
  END la_oenb[66]
  PIN la_oenb[67]
    PORT
      LAYER met2 ;
        RECT 1100.410 3296.000 1100.690 3300.000 ;
    END
  END la_oenb[67]
  PIN la_oenb[68]
    PORT
      LAYER met2 ;
        RECT 1115.590 3296.000 1115.870 3300.000 ;
    END
  END la_oenb[68]
  PIN la_oenb[69]
    PORT
      LAYER met2 ;
        RECT 1130.770 3296.000 1131.050 3300.000 ;
    END
  END la_oenb[69]
  PIN la_oenb[6]
    PORT
      LAYER met2 ;
        RECT 174.430 3296.000 174.710 3300.000 ;
    END
  END la_oenb[6]
  PIN la_oenb[70]
    PORT
      LAYER met2 ;
        RECT 1145.950 3296.000 1146.230 3300.000 ;
    END
  END la_oenb[70]
  PIN la_oenb[71]
    PORT
      LAYER met2 ;
        RECT 1161.130 3296.000 1161.410 3300.000 ;
    END
  END la_oenb[71]
  PIN la_oenb[72]
    PORT
      LAYER met2 ;
        RECT 1176.310 3296.000 1176.590 3300.000 ;
    END
  END la_oenb[72]
  PIN la_oenb[73]
    PORT
      LAYER met2 ;
        RECT 1191.490 3296.000 1191.770 3300.000 ;
    END
  END la_oenb[73]
  PIN la_oenb[74]
    PORT
      LAYER met2 ;
        RECT 1206.670 3296.000 1206.950 3300.000 ;
    END
  END la_oenb[74]
  PIN la_oenb[75]
    PORT
      LAYER met2 ;
        RECT 1221.850 3296.000 1222.130 3300.000 ;
    END
  END la_oenb[75]
  PIN la_oenb[76]
    PORT
      LAYER met2 ;
        RECT 1237.030 3296.000 1237.310 3300.000 ;
    END
  END la_oenb[76]
  PIN la_oenb[77]
    PORT
      LAYER met2 ;
        RECT 1252.210 3296.000 1252.490 3300.000 ;
    END
  END la_oenb[77]
  PIN la_oenb[78]
    PORT
      LAYER met2 ;
        RECT 1267.390 3296.000 1267.670 3300.000 ;
    END
  END la_oenb[78]
  PIN la_oenb[79]
    PORT
      LAYER met2 ;
        RECT 1282.570 3296.000 1282.850 3300.000 ;
    END
  END la_oenb[79]
  PIN la_oenb[7]
    PORT
      LAYER met2 ;
        RECT 189.610 3296.000 189.890 3300.000 ;
    END
  END la_oenb[7]
  PIN la_oenb[80]
    PORT
      LAYER met2 ;
        RECT 1297.750 3296.000 1298.030 3300.000 ;
    END
  END la_oenb[80]
  PIN la_oenb[81]
    PORT
      LAYER met2 ;
        RECT 1312.930 3296.000 1313.210 3300.000 ;
    END
  END la_oenb[81]
  PIN la_oenb[82]
    PORT
      LAYER met2 ;
        RECT 1328.110 3296.000 1328.390 3300.000 ;
    END
  END la_oenb[82]
  PIN la_oenb[83]
    PORT
      LAYER met2 ;
        RECT 1343.290 3296.000 1343.570 3300.000 ;
    END
  END la_oenb[83]
  PIN la_oenb[84]
    PORT
      LAYER met2 ;
        RECT 1358.470 3296.000 1358.750 3300.000 ;
    END
  END la_oenb[84]
  PIN la_oenb[85]
    PORT
      LAYER met2 ;
        RECT 1373.650 3296.000 1373.930 3300.000 ;
    END
  END la_oenb[85]
  PIN la_oenb[86]
    PORT
      LAYER met2 ;
        RECT 1388.830 3296.000 1389.110 3300.000 ;
    END
  END la_oenb[86]
  PIN la_oenb[87]
    PORT
      LAYER met2 ;
        RECT 1404.010 3296.000 1404.290 3300.000 ;
    END
  END la_oenb[87]
  PIN la_oenb[88]
    PORT
      LAYER met2 ;
        RECT 1419.190 3296.000 1419.470 3300.000 ;
    END
  END la_oenb[88]
  PIN la_oenb[89]
    PORT
      LAYER met2 ;
        RECT 1434.370 3296.000 1434.650 3300.000 ;
    END
  END la_oenb[89]
  PIN la_oenb[8]
    PORT
      LAYER met2 ;
        RECT 204.790 3296.000 205.070 3300.000 ;
    END
  END la_oenb[8]
  PIN la_oenb[90]
    PORT
      LAYER met2 ;
        RECT 1449.550 3296.000 1449.830 3300.000 ;
    END
  END la_oenb[90]
  PIN la_oenb[91]
    PORT
      LAYER met2 ;
        RECT 1464.730 3296.000 1465.010 3300.000 ;
    END
  END la_oenb[91]
  PIN la_oenb[92]
    PORT
      LAYER met2 ;
        RECT 1479.910 3296.000 1480.190 3300.000 ;
    END
  END la_oenb[92]
  PIN la_oenb[93]
    PORT
      LAYER met2 ;
        RECT 1495.090 3296.000 1495.370 3300.000 ;
    END
  END la_oenb[93]
  PIN la_oenb[94]
    PORT
      LAYER met2 ;
        RECT 1510.270 3296.000 1510.550 3300.000 ;
    END
  END la_oenb[94]
  PIN la_oenb[95]
    PORT
      LAYER met2 ;
        RECT 1525.450 3296.000 1525.730 3300.000 ;
    END
  END la_oenb[95]
  PIN la_oenb[96]
    PORT
      LAYER met2 ;
        RECT 1540.630 3296.000 1540.910 3300.000 ;
    END
  END la_oenb[96]
  PIN la_oenb[97]
    PORT
      LAYER met2 ;
        RECT 1555.810 3296.000 1556.090 3300.000 ;
    END
  END la_oenb[97]
  PIN la_oenb[98]
    PORT
      LAYER met2 ;
        RECT 1570.990 3296.000 1571.270 3300.000 ;
    END
  END la_oenb[98]
  PIN la_oenb[99]
    PORT
      LAYER met2 ;
        RECT 1586.170 3296.000 1586.450 3300.000 ;
    END
  END la_oenb[99]
  PIN la_oenb[9]
    PORT
      LAYER met2 ;
        RECT 219.970 3296.000 220.250 3300.000 ;
    END
  END la_oenb[9]
  PIN vccd1
    PORT
      LAYER met5 ;
        RECT 5.280 2822.080 2094.620 2823.680 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 3272.080 2094.620 3273.680 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 3197.080 2094.620 3198.680 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 3122.080 2094.620 3123.680 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 3047.080 2094.620 3048.680 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 2972.080 2094.620 2973.680 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 2897.080 2094.620 2898.680 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 2747.080 2094.620 2748.680 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 2672.080 2094.620 2673.680 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 2597.080 2094.620 2598.680 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 2522.080 2094.620 2523.680 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 2447.080 2094.620 2448.680 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 2372.080 2094.620 2373.680 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 2297.080 2094.620 2298.680 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 2222.080 2094.620 2223.680 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 2147.080 2094.620 2148.680 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 2072.080 2094.620 2073.680 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 1997.080 2094.620 1998.680 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 1922.080 2094.620 1923.680 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 1847.080 2094.620 1848.680 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 1772.080 2094.620 1773.680 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 1697.080 2094.620 1698.680 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 1622.080 2094.620 1623.680 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 1547.080 2094.620 1548.680 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 1472.080 2094.620 1473.680 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 1397.080 2094.620 1398.680 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 1322.080 2094.620 1323.680 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 1247.080 2094.620 1248.680 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 1172.080 2094.620 1173.680 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 1097.080 2094.620 1098.680 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 1022.080 2094.620 1023.680 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 947.080 2094.620 948.680 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 872.080 2094.620 873.680 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 797.080 2094.620 798.680 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 722.080 2094.620 723.680 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 647.080 2094.620 648.680 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 572.080 2094.620 573.680 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 497.080 2094.620 498.680 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 422.080 2094.620 423.680 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 347.080 2094.620 348.680 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 272.080 2094.620 273.680 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 197.080 2094.620 198.680 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 122.080 2094.620 123.680 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 47.080 2094.620 48.680 ;
    END
    PORT
      LAYER met4 ;
        RECT 2071.720 10.640 2073.320 3288.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 2001.720 10.640 2003.320 3288.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 1931.720 10.640 1933.320 3288.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 1861.720 2887.580 1863.320 3288.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 1861.720 2687.580 1863.320 2810.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 1861.720 2487.580 1863.320 2610.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 1861.720 2287.580 1863.320 2410.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 1861.720 2087.580 1863.320 2210.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 1861.720 1887.580 1863.320 2010.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 1861.720 1687.580 1863.320 1810.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 1861.720 1487.580 1863.320 1610.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 1861.720 1287.580 1863.320 1410.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 1861.720 1087.580 1863.320 1210.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 1861.720 887.580 1863.320 1010.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 1861.720 687.580 1863.320 810.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 1861.720 487.580 1863.320 610.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 1861.720 10.640 1863.320 410.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 1791.720 10.640 1793.320 3288.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 1721.720 10.640 1723.320 3288.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 1651.720 2890.185 1653.320 3288.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 1651.720 2277.265 1653.320 2836.295 ;
    END
    PORT
      LAYER met4 ;
        RECT 1651.720 1677.265 1653.320 2230.175 ;
    END
    PORT
      LAYER met4 ;
        RECT 1651.720 1077.265 1653.320 1630.175 ;
    END
    PORT
      LAYER met4 ;
        RECT 1651.720 10.640 1653.320 1030.175 ;
    END
    PORT
      LAYER met4 ;
        RECT 1581.720 10.640 1583.320 3288.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 1511.720 10.640 1513.320 3288.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 1441.720 2684.065 1443.320 3288.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 1441.720 2284.065 1443.320 2611.815 ;
    END
    PORT
      LAYER met4 ;
        RECT 1441.720 2084.065 1443.320 2205.695 ;
    END
    PORT
      LAYER met4 ;
        RECT 1441.720 1684.065 1443.320 2011.815 ;
    END
    PORT
      LAYER met4 ;
        RECT 1441.720 1484.065 1443.320 1605.695 ;
    END
    PORT
      LAYER met4 ;
        RECT 1441.720 1084.065 1443.320 1411.815 ;
    END
    PORT
      LAYER met4 ;
        RECT 1441.720 884.065 1443.320 1005.695 ;
    END
    PORT
      LAYER met4 ;
        RECT 1441.720 10.640 1443.320 811.815 ;
    END
    PORT
      LAYER met4 ;
        RECT 1371.720 10.640 1373.320 3288.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 1301.720 2698.460 1303.320 3288.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 1301.720 2098.460 1303.320 2610.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 1301.720 1498.460 1303.320 2010.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 1301.720 898.460 1303.320 1410.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 1301.720 10.640 1303.320 810.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 1231.720 2890.185 1233.320 3288.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 1231.720 2277.265 1233.320 2836.295 ;
    END
    PORT
      LAYER met4 ;
        RECT 1231.720 1677.265 1233.320 2230.175 ;
    END
    PORT
      LAYER met4 ;
        RECT 1231.720 1077.265 1233.320 1630.175 ;
    END
    PORT
      LAYER met4 ;
        RECT 1231.720 10.640 1233.320 1030.175 ;
    END
    PORT
      LAYER met4 ;
        RECT 1161.720 10.640 1163.320 3288.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 1091.720 2887.580 1093.320 3288.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 1091.720 2687.580 1093.320 2810.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 1091.720 2287.580 1093.320 2610.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 1091.720 2087.580 1093.320 2205.695 ;
    END
    PORT
      LAYER met4 ;
        RECT 1091.720 1687.580 1093.320 2010.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 1091.720 1487.580 1093.320 1605.695 ;
    END
    PORT
      LAYER met4 ;
        RECT 1091.720 1087.580 1093.320 1410.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 1091.720 887.580 1093.320 1005.695 ;
    END
    PORT
      LAYER met4 ;
        RECT 1091.720 487.580 1093.320 810.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 1091.720 10.640 1093.320 410.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 1021.720 2684.065 1023.320 3288.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 1021.720 2284.065 1023.320 2611.815 ;
    END
    PORT
      LAYER met4 ;
        RECT 1021.720 2084.065 1023.320 2205.695 ;
    END
    PORT
      LAYER met4 ;
        RECT 1021.720 1684.065 1023.320 2011.815 ;
    END
    PORT
      LAYER met4 ;
        RECT 1021.720 1484.065 1023.320 1605.695 ;
    END
    PORT
      LAYER met4 ;
        RECT 1021.720 1084.065 1023.320 1411.815 ;
    END
    PORT
      LAYER met4 ;
        RECT 1021.720 884.065 1023.320 1005.695 ;
    END
    PORT
      LAYER met4 ;
        RECT 1021.720 10.640 1023.320 811.815 ;
    END
    PORT
      LAYER met4 ;
        RECT 951.720 10.640 953.320 3288.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 881.720 3087.580 883.320 3288.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 881.720 2890.185 883.320 3010.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 881.720 2687.465 883.320 2810.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 881.720 2287.580 883.320 2616.575 ;
    END
    PORT
      LAYER met4 ;
        RECT 881.720 2087.465 883.320 2210.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 881.720 1687.580 883.320 2016.575 ;
    END
    PORT
      LAYER met4 ;
        RECT 881.720 1487.465 883.320 1610.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 881.720 1087.580 883.320 1416.575 ;
    END
    PORT
      LAYER met4 ;
        RECT 881.720 887.465 883.320 1010.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 881.720 487.580 883.320 816.575 ;
    END
    PORT
      LAYER met4 ;
        RECT 881.720 287.580 883.320 410.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 881.720 10.640 883.320 210.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 811.720 2890.185 813.320 3288.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 811.720 10.640 813.320 2836.295 ;
    END
    PORT
      LAYER met4 ;
        RECT 741.720 10.640 743.320 3288.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 671.720 2887.580 673.320 3288.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 671.720 2687.580 673.320 2810.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 671.720 2287.580 673.320 2610.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 671.720 2087.580 673.320 2205.695 ;
    END
    PORT
      LAYER met4 ;
        RECT 671.720 1687.580 673.320 2010.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 671.720 1487.580 673.320 1605.695 ;
    END
    PORT
      LAYER met4 ;
        RECT 671.720 1087.580 673.320 1410.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 671.720 887.580 673.320 1005.695 ;
    END
    PORT
      LAYER met4 ;
        RECT 671.720 487.580 673.320 810.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 671.720 10.640 673.320 410.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 601.720 10.640 603.320 3288.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 531.720 10.640 533.320 3288.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 461.720 3087.580 463.320 3288.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 461.720 2890.185 463.320 3010.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 461.720 2287.580 463.320 2810.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 461.720 1687.580 463.320 2210.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 461.720 1087.580 463.320 1610.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 461.720 487.580 463.320 1010.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 461.720 287.580 463.320 410.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 461.720 10.640 463.320 210.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 391.720 10.640 393.320 3288.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 321.720 10.640 323.320 3288.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.720 10.640 253.320 3288.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 181.720 10.640 183.320 3288.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 111.720 10.640 113.320 3288.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 41.720 10.640 43.320 3288.720 ;
    END
  END vccd1
  PIN vssd1
    PORT
      LAYER met5 ;
        RECT 5.280 2825.380 2094.620 2826.980 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 3275.380 2094.620 3276.980 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 3200.380 2094.620 3201.980 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 3125.380 2094.620 3126.980 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 3050.380 2094.620 3051.980 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 2975.380 2094.620 2976.980 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 2900.380 2094.620 2901.980 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 2750.380 2094.620 2751.980 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 2675.380 2094.620 2676.980 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 2600.380 2094.620 2601.980 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 2525.380 2094.620 2526.980 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 2450.380 2094.620 2451.980 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 2375.380 2094.620 2376.980 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 2300.380 2094.620 2301.980 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 2225.380 2094.620 2226.980 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 2150.380 2094.620 2151.980 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 2075.380 2094.620 2076.980 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 2000.380 2094.620 2001.980 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 1925.380 2094.620 1926.980 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 1850.380 2094.620 1851.980 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 1775.380 2094.620 1776.980 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 1700.380 2094.620 1701.980 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 1625.380 2094.620 1626.980 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 1550.380 2094.620 1551.980 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 1475.380 2094.620 1476.980 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 1400.380 2094.620 1401.980 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 1325.380 2094.620 1326.980 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 1250.380 2094.620 1251.980 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 1175.380 2094.620 1176.980 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 1100.380 2094.620 1101.980 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 1025.380 2094.620 1026.980 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 950.380 2094.620 951.980 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 875.380 2094.620 876.980 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 800.380 2094.620 801.980 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 725.380 2094.620 726.980 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 650.380 2094.620 651.980 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 575.380 2094.620 576.980 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 500.380 2094.620 501.980 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 425.380 2094.620 426.980 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 350.380 2094.620 351.980 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 275.380 2094.620 276.980 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 200.380 2094.620 201.980 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 125.380 2094.620 126.980 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 50.380 2094.620 51.980 ;
    END
    PORT
      LAYER met4 ;
        RECT 2075.020 10.640 2076.620 3288.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 2005.020 10.640 2006.620 3288.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 1935.020 10.640 1936.620 3288.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 1865.020 2849.385 1866.620 3288.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 1865.020 2684.065 1866.620 2826.095 ;
    END
    PORT
      LAYER met4 ;
        RECT 1865.020 2084.065 1866.620 2611.815 ;
    END
    PORT
      LAYER met4 ;
        RECT 1865.020 1484.065 1866.620 2011.815 ;
    END
    PORT
      LAYER met4 ;
        RECT 1865.020 884.065 1866.620 1411.815 ;
    END
    PORT
      LAYER met4 ;
        RECT 1865.020 10.640 1866.620 811.815 ;
    END
    PORT
      LAYER met4 ;
        RECT 1795.020 10.640 1796.620 3288.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 1725.020 10.640 1726.620 3288.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 1655.020 2890.185 1656.620 3288.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 1655.020 2698.460 1656.620 2836.295 ;
    END
    PORT
      LAYER met4 ;
        RECT 1655.020 2277.265 1656.620 2610.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 1655.020 2098.460 1656.620 2230.175 ;
    END
    PORT
      LAYER met4 ;
        RECT 1655.020 1677.265 1656.620 2010.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 1655.020 1498.460 1656.620 1630.175 ;
    END
    PORT
      LAYER met4 ;
        RECT 1655.020 1077.265 1656.620 1410.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 1655.020 898.460 1656.620 1030.175 ;
    END
    PORT
      LAYER met4 ;
        RECT 1655.020 10.640 1656.620 810.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 1585.020 10.640 1586.620 3288.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 1515.020 10.640 1516.620 3288.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 1445.020 2684.065 1446.620 3288.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 1445.020 2284.065 1446.620 2611.815 ;
    END
    PORT
      LAYER met4 ;
        RECT 1445.020 2084.065 1446.620 2205.695 ;
    END
    PORT
      LAYER met4 ;
        RECT 1445.020 1684.065 1446.620 2011.815 ;
    END
    PORT
      LAYER met4 ;
        RECT 1445.020 1484.065 1446.620 1605.695 ;
    END
    PORT
      LAYER met4 ;
        RECT 1445.020 1084.065 1446.620 1411.815 ;
    END
    PORT
      LAYER met4 ;
        RECT 1445.020 884.065 1446.620 1005.695 ;
    END
    PORT
      LAYER met4 ;
        RECT 1445.020 10.640 1446.620 811.815 ;
    END
    PORT
      LAYER met4 ;
        RECT 1375.020 10.640 1376.620 3288.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 1305.020 2698.460 1306.620 3288.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 1305.020 2098.460 1306.620 2610.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 1305.020 1498.460 1306.620 2010.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 1305.020 898.460 1306.620 1410.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 1305.020 10.640 1306.620 810.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 1235.020 2890.185 1236.620 3288.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 1235.020 2277.265 1236.620 2836.295 ;
    END
    PORT
      LAYER met4 ;
        RECT 1235.020 1677.265 1236.620 2230.175 ;
    END
    PORT
      LAYER met4 ;
        RECT 1235.020 1077.265 1236.620 1630.175 ;
    END
    PORT
      LAYER met4 ;
        RECT 1235.020 10.640 1236.620 1030.175 ;
    END
    PORT
      LAYER met4 ;
        RECT 1165.020 10.640 1166.620 3288.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 1095.020 2887.580 1096.620 3288.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 1095.020 2687.580 1096.620 2810.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 1095.020 2287.580 1096.620 2610.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 1095.020 2087.580 1096.620 2205.695 ;
    END
    PORT
      LAYER met4 ;
        RECT 1095.020 1687.580 1096.620 2010.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 1095.020 1487.580 1096.620 1605.695 ;
    END
    PORT
      LAYER met4 ;
        RECT 1095.020 1087.580 1096.620 1410.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 1095.020 887.580 1096.620 1005.695 ;
    END
    PORT
      LAYER met4 ;
        RECT 1095.020 487.580 1096.620 810.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 1095.020 10.640 1096.620 410.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 1025.020 2887.580 1026.620 3288.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 1025.020 2687.580 1026.620 2810.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 1025.020 2287.580 1026.620 2610.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 1025.020 2087.580 1026.620 2205.695 ;
    END
    PORT
      LAYER met4 ;
        RECT 1025.020 1687.580 1026.620 2010.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 1025.020 1487.580 1026.620 1605.695 ;
    END
    PORT
      LAYER met4 ;
        RECT 1025.020 1087.580 1026.620 1410.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 1025.020 887.580 1026.620 1005.695 ;
    END
    PORT
      LAYER met4 ;
        RECT 1025.020 487.580 1026.620 810.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 1025.020 10.640 1026.620 410.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 955.020 10.640 956.620 3288.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 885.020 2890.185 886.620 3288.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 885.020 2687.465 886.620 2836.295 ;
    END
    PORT
      LAYER met4 ;
        RECT 885.020 2087.465 886.620 2616.575 ;
    END
    PORT
      LAYER met4 ;
        RECT 885.020 1487.465 886.620 2016.575 ;
    END
    PORT
      LAYER met4 ;
        RECT 885.020 887.465 886.620 1416.575 ;
    END
    PORT
      LAYER met4 ;
        RECT 885.020 437.145 886.620 816.575 ;
    END
    PORT
      LAYER met4 ;
        RECT 885.020 10.640 886.620 426.775 ;
    END
    PORT
      LAYER met4 ;
        RECT 815.020 3087.580 816.620 3288.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 815.020 2890.185 816.620 3010.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 815.020 2698.460 816.620 2810.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 815.020 2287.580 816.620 2610.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 815.020 2098.460 816.620 2210.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 815.020 1687.580 816.620 2010.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 815.020 1498.460 816.620 1610.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 815.020 1087.580 816.620 1410.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 815.020 898.460 816.620 1010.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 815.020 487.580 816.620 810.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 815.020 287.580 816.620 410.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 815.020 10.640 816.620 210.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 745.020 10.640 746.620 3288.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 675.020 2880.665 676.620 3288.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 675.020 2684.065 676.620 2812.495 ;
    END
    PORT
      LAYER met4 ;
        RECT 675.020 2284.065 676.620 2611.815 ;
    END
    PORT
      LAYER met4 ;
        RECT 675.020 2084.065 676.620 2205.695 ;
    END
    PORT
      LAYER met4 ;
        RECT 675.020 1684.065 676.620 2011.815 ;
    END
    PORT
      LAYER met4 ;
        RECT 675.020 1484.065 676.620 1605.695 ;
    END
    PORT
      LAYER met4 ;
        RECT 675.020 1084.065 676.620 1411.815 ;
    END
    PORT
      LAYER met4 ;
        RECT 675.020 884.065 676.620 1005.695 ;
    END
    PORT
      LAYER met4 ;
        RECT 675.020 471.825 676.620 811.815 ;
    END
    PORT
      LAYER met4 ;
        RECT 675.020 10.640 676.620 427.455 ;
    END
    PORT
      LAYER met4 ;
        RECT 605.020 2684.065 606.620 3288.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 605.020 2284.065 606.620 2611.815 ;
    END
    PORT
      LAYER met4 ;
        RECT 605.020 2084.065 606.620 2205.695 ;
    END
    PORT
      LAYER met4 ;
        RECT 605.020 1684.065 606.620 2011.815 ;
    END
    PORT
      LAYER met4 ;
        RECT 605.020 1484.065 606.620 1605.695 ;
    END
    PORT
      LAYER met4 ;
        RECT 605.020 1084.065 606.620 1411.815 ;
    END
    PORT
      LAYER met4 ;
        RECT 605.020 884.065 606.620 1005.695 ;
    END
    PORT
      LAYER met4 ;
        RECT 605.020 10.640 606.620 811.815 ;
    END
    PORT
      LAYER met4 ;
        RECT 535.020 10.640 536.620 3288.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 465.020 2890.185 466.620 3288.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 465.020 2698.460 466.620 2836.295 ;
    END
    PORT
      LAYER met4 ;
        RECT 465.020 2098.460 466.620 2610.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 465.020 1498.460 466.620 2010.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 465.020 898.460 466.620 1410.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 465.020 10.640 466.620 810.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 395.020 10.640 396.620 3288.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 325.020 10.640 326.620 3288.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 255.020 10.640 256.620 3288.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 185.020 10.640 186.620 3288.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 115.020 10.640 116.620 3288.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 45.020 10.640 46.620 3288.720 ;
    END
  END vssd1
  PIN wb_clk_i
    PORT
      LAYER met2 ;
        RECT 11.130 0.000 11.410 4.000 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    PORT
      LAYER met2 ;
        RECT 30.910 0.000 31.190 4.000 ;
    END
  END wb_rst_i
  PIN wbs_ack_o
    PORT
      LAYER met2 ;
        RECT 50.690 0.000 50.970 4.000 ;
    END
  END wbs_ack_o
  PIN wbs_adr_i[0]
    PORT
      LAYER met2 ;
        RECT 129.810 0.000 130.090 4.000 ;
    END
  END wbs_adr_i[0]
  PIN wbs_adr_i[10]
    PORT
      LAYER met2 ;
        RECT 802.330 0.000 802.610 4.000 ;
    END
  END wbs_adr_i[10]
  PIN wbs_adr_i[11]
    PORT
      LAYER met2 ;
        RECT 861.670 0.000 861.950 4.000 ;
    END
  END wbs_adr_i[11]
  PIN wbs_adr_i[12]
    PORT
      LAYER met2 ;
        RECT 921.010 0.000 921.290 4.000 ;
    END
  END wbs_adr_i[12]
  PIN wbs_adr_i[13]
    PORT
      LAYER met2 ;
        RECT 980.350 0.000 980.630 4.000 ;
    END
  END wbs_adr_i[13]
  PIN wbs_adr_i[14]
    PORT
      LAYER met2 ;
        RECT 1039.690 0.000 1039.970 4.000 ;
    END
  END wbs_adr_i[14]
  PIN wbs_adr_i[15]
    PORT
      LAYER met2 ;
        RECT 1099.030 0.000 1099.310 4.000 ;
    END
  END wbs_adr_i[15]
  PIN wbs_adr_i[16]
    PORT
      LAYER met2 ;
        RECT 1158.370 0.000 1158.650 4.000 ;
    END
  END wbs_adr_i[16]
  PIN wbs_adr_i[17]
    PORT
      LAYER met2 ;
        RECT 1217.710 0.000 1217.990 4.000 ;
    END
  END wbs_adr_i[17]
  PIN wbs_adr_i[18]
    PORT
      LAYER met2 ;
        RECT 1277.050 0.000 1277.330 4.000 ;
    END
  END wbs_adr_i[18]
  PIN wbs_adr_i[19]
    PORT
      LAYER met2 ;
        RECT 1336.390 0.000 1336.670 4.000 ;
    END
  END wbs_adr_i[19]
  PIN wbs_adr_i[1]
    PORT
      LAYER met2 ;
        RECT 208.930 0.000 209.210 4.000 ;
    END
  END wbs_adr_i[1]
  PIN wbs_adr_i[20]
    PORT
      LAYER met2 ;
        RECT 1395.730 0.000 1396.010 4.000 ;
    END
  END wbs_adr_i[20]
  PIN wbs_adr_i[21]
    PORT
      LAYER met2 ;
        RECT 1455.070 0.000 1455.350 4.000 ;
    END
  END wbs_adr_i[21]
  PIN wbs_adr_i[22]
    PORT
      LAYER met2 ;
        RECT 1514.410 0.000 1514.690 4.000 ;
    END
  END wbs_adr_i[22]
  PIN wbs_adr_i[23]
    PORT
      LAYER met2 ;
        RECT 1573.750 0.000 1574.030 4.000 ;
    END
  END wbs_adr_i[23]
  PIN wbs_adr_i[24]
    PORT
      LAYER met2 ;
        RECT 1633.090 0.000 1633.370 4.000 ;
    END
  END wbs_adr_i[24]
  PIN wbs_adr_i[25]
    PORT
      LAYER met2 ;
        RECT 1692.430 0.000 1692.710 4.000 ;
    END
  END wbs_adr_i[25]
  PIN wbs_adr_i[26]
    PORT
      LAYER met2 ;
        RECT 1751.770 0.000 1752.050 4.000 ;
    END
  END wbs_adr_i[26]
  PIN wbs_adr_i[27]
    PORT
      LAYER met2 ;
        RECT 1811.110 0.000 1811.390 4.000 ;
    END
  END wbs_adr_i[27]
  PIN wbs_adr_i[28]
    PORT
      LAYER met2 ;
        RECT 1870.450 0.000 1870.730 4.000 ;
    END
  END wbs_adr_i[28]
  PIN wbs_adr_i[29]
    PORT
      LAYER met2 ;
        RECT 1929.790 0.000 1930.070 4.000 ;
    END
  END wbs_adr_i[29]
  PIN wbs_adr_i[2]
    PORT
      LAYER met2 ;
        RECT 288.050 0.000 288.330 4.000 ;
    END
  END wbs_adr_i[2]
  PIN wbs_adr_i[30]
    PORT
      LAYER met2 ;
        RECT 1989.130 0.000 1989.410 4.000 ;
    END
  END wbs_adr_i[30]
  PIN wbs_adr_i[31]
    PORT
      LAYER met2 ;
        RECT 2048.470 0.000 2048.750 4.000 ;
    END
  END wbs_adr_i[31]
  PIN wbs_adr_i[3]
    PORT
      LAYER met2 ;
        RECT 367.170 0.000 367.450 4.000 ;
    END
  END wbs_adr_i[3]
  PIN wbs_adr_i[4]
    PORT
      LAYER met2 ;
        RECT 446.290 0.000 446.570 4.000 ;
    END
  END wbs_adr_i[4]
  PIN wbs_adr_i[5]
    PORT
      LAYER met2 ;
        RECT 505.630 0.000 505.910 4.000 ;
    END
  END wbs_adr_i[5]
  PIN wbs_adr_i[6]
    PORT
      LAYER met2 ;
        RECT 564.970 0.000 565.250 4.000 ;
    END
  END wbs_adr_i[6]
  PIN wbs_adr_i[7]
    PORT
      LAYER met2 ;
        RECT 624.310 0.000 624.590 4.000 ;
    END
  END wbs_adr_i[7]
  PIN wbs_adr_i[8]
    PORT
      LAYER met2 ;
        RECT 683.650 0.000 683.930 4.000 ;
    END
  END wbs_adr_i[8]
  PIN wbs_adr_i[9]
    PORT
      LAYER met2 ;
        RECT 742.990 0.000 743.270 4.000 ;
    END
  END wbs_adr_i[9]
  PIN wbs_cyc_i
    PORT
      LAYER met2 ;
        RECT 70.470 0.000 70.750 4.000 ;
    END
  END wbs_cyc_i
  PIN wbs_dat_i[0]
    PORT
      LAYER met2 ;
        RECT 149.590 0.000 149.870 4.000 ;
    END
  END wbs_dat_i[0]
  PIN wbs_dat_i[10]
    PORT
      LAYER met2 ;
        RECT 822.110 0.000 822.390 4.000 ;
    END
  END wbs_dat_i[10]
  PIN wbs_dat_i[11]
    PORT
      LAYER met2 ;
        RECT 881.450 0.000 881.730 4.000 ;
    END
  END wbs_dat_i[11]
  PIN wbs_dat_i[12]
    PORT
      LAYER met2 ;
        RECT 940.790 0.000 941.070 4.000 ;
    END
  END wbs_dat_i[12]
  PIN wbs_dat_i[13]
    PORT
      LAYER met2 ;
        RECT 1000.130 0.000 1000.410 4.000 ;
    END
  END wbs_dat_i[13]
  PIN wbs_dat_i[14]
    PORT
      LAYER met2 ;
        RECT 1059.470 0.000 1059.750 4.000 ;
    END
  END wbs_dat_i[14]
  PIN wbs_dat_i[15]
    PORT
      LAYER met2 ;
        RECT 1118.810 0.000 1119.090 4.000 ;
    END
  END wbs_dat_i[15]
  PIN wbs_dat_i[16]
    PORT
      LAYER met2 ;
        RECT 1178.150 0.000 1178.430 4.000 ;
    END
  END wbs_dat_i[16]
  PIN wbs_dat_i[17]
    PORT
      LAYER met2 ;
        RECT 1237.490 0.000 1237.770 4.000 ;
    END
  END wbs_dat_i[17]
  PIN wbs_dat_i[18]
    PORT
      LAYER met2 ;
        RECT 1296.830 0.000 1297.110 4.000 ;
    END
  END wbs_dat_i[18]
  PIN wbs_dat_i[19]
    PORT
      LAYER met2 ;
        RECT 1356.170 0.000 1356.450 4.000 ;
    END
  END wbs_dat_i[19]
  PIN wbs_dat_i[1]
    PORT
      LAYER met2 ;
        RECT 228.710 0.000 228.990 4.000 ;
    END
  END wbs_dat_i[1]
  PIN wbs_dat_i[20]
    PORT
      LAYER met2 ;
        RECT 1415.510 0.000 1415.790 4.000 ;
    END
  END wbs_dat_i[20]
  PIN wbs_dat_i[21]
    PORT
      LAYER met2 ;
        RECT 1474.850 0.000 1475.130 4.000 ;
    END
  END wbs_dat_i[21]
  PIN wbs_dat_i[22]
    PORT
      LAYER met2 ;
        RECT 1534.190 0.000 1534.470 4.000 ;
    END
  END wbs_dat_i[22]
  PIN wbs_dat_i[23]
    PORT
      LAYER met2 ;
        RECT 1593.530 0.000 1593.810 4.000 ;
    END
  END wbs_dat_i[23]
  PIN wbs_dat_i[24]
    PORT
      LAYER met2 ;
        RECT 1652.870 0.000 1653.150 4.000 ;
    END
  END wbs_dat_i[24]
  PIN wbs_dat_i[25]
    PORT
      LAYER met2 ;
        RECT 1712.210 0.000 1712.490 4.000 ;
    END
  END wbs_dat_i[25]
  PIN wbs_dat_i[26]
    PORT
      LAYER met2 ;
        RECT 1771.550 0.000 1771.830 4.000 ;
    END
  END wbs_dat_i[26]
  PIN wbs_dat_i[27]
    PORT
      LAYER met2 ;
        RECT 1830.890 0.000 1831.170 4.000 ;
    END
  END wbs_dat_i[27]
  PIN wbs_dat_i[28]
    PORT
      LAYER met2 ;
        RECT 1890.230 0.000 1890.510 4.000 ;
    END
  END wbs_dat_i[28]
  PIN wbs_dat_i[29]
    PORT
      LAYER met2 ;
        RECT 1949.570 0.000 1949.850 4.000 ;
    END
  END wbs_dat_i[29]
  PIN wbs_dat_i[2]
    PORT
      LAYER met2 ;
        RECT 307.830 0.000 308.110 4.000 ;
    END
  END wbs_dat_i[2]
  PIN wbs_dat_i[30]
    PORT
      LAYER met2 ;
        RECT 2008.910 0.000 2009.190 4.000 ;
    END
  END wbs_dat_i[30]
  PIN wbs_dat_i[31]
    PORT
      LAYER met2 ;
        RECT 2068.250 0.000 2068.530 4.000 ;
    END
  END wbs_dat_i[31]
  PIN wbs_dat_i[3]
    PORT
      LAYER met2 ;
        RECT 386.950 0.000 387.230 4.000 ;
    END
  END wbs_dat_i[3]
  PIN wbs_dat_i[4]
    PORT
      LAYER met2 ;
        RECT 466.070 0.000 466.350 4.000 ;
    END
  END wbs_dat_i[4]
  PIN wbs_dat_i[5]
    PORT
      LAYER met2 ;
        RECT 525.410 0.000 525.690 4.000 ;
    END
  END wbs_dat_i[5]
  PIN wbs_dat_i[6]
    PORT
      LAYER met2 ;
        RECT 584.750 0.000 585.030 4.000 ;
    END
  END wbs_dat_i[6]
  PIN wbs_dat_i[7]
    PORT
      LAYER met2 ;
        RECT 644.090 0.000 644.370 4.000 ;
    END
  END wbs_dat_i[7]
  PIN wbs_dat_i[8]
    PORT
      LAYER met2 ;
        RECT 703.430 0.000 703.710 4.000 ;
    END
  END wbs_dat_i[8]
  PIN wbs_dat_i[9]
    PORT
      LAYER met2 ;
        RECT 762.770 0.000 763.050 4.000 ;
    END
  END wbs_dat_i[9]
  PIN wbs_dat_o[0]
    PORT
      LAYER met2 ;
        RECT 169.370 0.000 169.650 4.000 ;
    END
  END wbs_dat_o[0]
  PIN wbs_dat_o[10]
    PORT
      LAYER met2 ;
        RECT 841.890 0.000 842.170 4.000 ;
    END
  END wbs_dat_o[10]
  PIN wbs_dat_o[11]
    PORT
      LAYER met2 ;
        RECT 901.230 0.000 901.510 4.000 ;
    END
  END wbs_dat_o[11]
  PIN wbs_dat_o[12]
    PORT
      LAYER met2 ;
        RECT 960.570 0.000 960.850 4.000 ;
    END
  END wbs_dat_o[12]
  PIN wbs_dat_o[13]
    PORT
      LAYER met2 ;
        RECT 1019.910 0.000 1020.190 4.000 ;
    END
  END wbs_dat_o[13]
  PIN wbs_dat_o[14]
    PORT
      LAYER met2 ;
        RECT 1079.250 0.000 1079.530 4.000 ;
    END
  END wbs_dat_o[14]
  PIN wbs_dat_o[15]
    PORT
      LAYER met2 ;
        RECT 1138.590 0.000 1138.870 4.000 ;
    END
  END wbs_dat_o[15]
  PIN wbs_dat_o[16]
    PORT
      LAYER met2 ;
        RECT 1197.930 0.000 1198.210 4.000 ;
    END
  END wbs_dat_o[16]
  PIN wbs_dat_o[17]
    PORT
      LAYER met2 ;
        RECT 1257.270 0.000 1257.550 4.000 ;
    END
  END wbs_dat_o[17]
  PIN wbs_dat_o[18]
    PORT
      LAYER met2 ;
        RECT 1316.610 0.000 1316.890 4.000 ;
    END
  END wbs_dat_o[18]
  PIN wbs_dat_o[19]
    PORT
      LAYER met2 ;
        RECT 1375.950 0.000 1376.230 4.000 ;
    END
  END wbs_dat_o[19]
  PIN wbs_dat_o[1]
    PORT
      LAYER met2 ;
        RECT 248.490 0.000 248.770 4.000 ;
    END
  END wbs_dat_o[1]
  PIN wbs_dat_o[20]
    PORT
      LAYER met2 ;
        RECT 1435.290 0.000 1435.570 4.000 ;
    END
  END wbs_dat_o[20]
  PIN wbs_dat_o[21]
    PORT
      LAYER met2 ;
        RECT 1494.630 0.000 1494.910 4.000 ;
    END
  END wbs_dat_o[21]
  PIN wbs_dat_o[22]
    PORT
      LAYER met2 ;
        RECT 1553.970 0.000 1554.250 4.000 ;
    END
  END wbs_dat_o[22]
  PIN wbs_dat_o[23]
    PORT
      LAYER met2 ;
        RECT 1613.310 0.000 1613.590 4.000 ;
    END
  END wbs_dat_o[23]
  PIN wbs_dat_o[24]
    PORT
      LAYER met2 ;
        RECT 1672.650 0.000 1672.930 4.000 ;
    END
  END wbs_dat_o[24]
  PIN wbs_dat_o[25]
    PORT
      LAYER met2 ;
        RECT 1731.990 0.000 1732.270 4.000 ;
    END
  END wbs_dat_o[25]
  PIN wbs_dat_o[26]
    PORT
      LAYER met2 ;
        RECT 1791.330 0.000 1791.610 4.000 ;
    END
  END wbs_dat_o[26]
  PIN wbs_dat_o[27]
    PORT
      LAYER met2 ;
        RECT 1850.670 0.000 1850.950 4.000 ;
    END
  END wbs_dat_o[27]
  PIN wbs_dat_o[28]
    PORT
      LAYER met2 ;
        RECT 1910.010 0.000 1910.290 4.000 ;
    END
  END wbs_dat_o[28]
  PIN wbs_dat_o[29]
    PORT
      LAYER met2 ;
        RECT 1969.350 0.000 1969.630 4.000 ;
    END
  END wbs_dat_o[29]
  PIN wbs_dat_o[2]
    PORT
      LAYER met2 ;
        RECT 327.610 0.000 327.890 4.000 ;
    END
  END wbs_dat_o[2]
  PIN wbs_dat_o[30]
    PORT
      LAYER met2 ;
        RECT 2028.690 0.000 2028.970 4.000 ;
    END
  END wbs_dat_o[30]
  PIN wbs_dat_o[31]
    PORT
      LAYER met2 ;
        RECT 2088.030 0.000 2088.310 4.000 ;
    END
  END wbs_dat_o[31]
  PIN wbs_dat_o[3]
    PORT
      LAYER met2 ;
        RECT 406.730 0.000 407.010 4.000 ;
    END
  END wbs_dat_o[3]
  PIN wbs_dat_o[4]
    PORT
      LAYER met2 ;
        RECT 485.850 0.000 486.130 4.000 ;
    END
  END wbs_dat_o[4]
  PIN wbs_dat_o[5]
    PORT
      LAYER met2 ;
        RECT 545.190 0.000 545.470 4.000 ;
    END
  END wbs_dat_o[5]
  PIN wbs_dat_o[6]
    PORT
      LAYER met2 ;
        RECT 604.530 0.000 604.810 4.000 ;
    END
  END wbs_dat_o[6]
  PIN wbs_dat_o[7]
    PORT
      LAYER met2 ;
        RECT 663.870 0.000 664.150 4.000 ;
    END
  END wbs_dat_o[7]
  PIN wbs_dat_o[8]
    PORT
      LAYER met2 ;
        RECT 723.210 0.000 723.490 4.000 ;
    END
  END wbs_dat_o[8]
  PIN wbs_dat_o[9]
    PORT
      LAYER met2 ;
        RECT 782.550 0.000 782.830 4.000 ;
    END
  END wbs_dat_o[9]
  PIN wbs_sel_i[0]
    PORT
      LAYER met2 ;
        RECT 189.150 0.000 189.430 4.000 ;
    END
  END wbs_sel_i[0]
  PIN wbs_sel_i[1]
    PORT
      LAYER met2 ;
        RECT 268.270 0.000 268.550 4.000 ;
    END
  END wbs_sel_i[1]
  PIN wbs_sel_i[2]
    PORT
      LAYER met2 ;
        RECT 347.390 0.000 347.670 4.000 ;
    END
  END wbs_sel_i[2]
  PIN wbs_sel_i[3]
    PORT
      LAYER met2 ;
        RECT 426.510 0.000 426.790 4.000 ;
    END
  END wbs_sel_i[3]
  PIN wbs_stb_i
    PORT
      LAYER met2 ;
        RECT 90.250 0.000 90.530 4.000 ;
    END
  END wbs_stb_i
  PIN wbs_we_i
    PORT
      LAYER met2 ;
        RECT 110.030 0.000 110.310 4.000 ;
    END
  END wbs_we_i
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 2094.380 3288.565 ;
      LAYER met1 ;
        RECT 4.670 10.640 2094.380 3288.720 ;
      LAYER met2 ;
        RECT 4.690 3295.720 72.950 3296.370 ;
        RECT 73.790 3295.720 78.010 3296.370 ;
        RECT 78.850 3295.720 83.070 3296.370 ;
        RECT 83.910 3295.720 88.130 3296.370 ;
        RECT 88.970 3295.720 93.190 3296.370 ;
        RECT 94.030 3295.720 98.250 3296.370 ;
        RECT 99.090 3295.720 103.310 3296.370 ;
        RECT 104.150 3295.720 108.370 3296.370 ;
        RECT 109.210 3295.720 113.430 3296.370 ;
        RECT 114.270 3295.720 118.490 3296.370 ;
        RECT 119.330 3295.720 123.550 3296.370 ;
        RECT 124.390 3295.720 128.610 3296.370 ;
        RECT 129.450 3295.720 133.670 3296.370 ;
        RECT 134.510 3295.720 138.730 3296.370 ;
        RECT 139.570 3295.720 143.790 3296.370 ;
        RECT 144.630 3295.720 148.850 3296.370 ;
        RECT 149.690 3295.720 153.910 3296.370 ;
        RECT 154.750 3295.720 158.970 3296.370 ;
        RECT 159.810 3295.720 164.030 3296.370 ;
        RECT 164.870 3295.720 169.090 3296.370 ;
        RECT 169.930 3295.720 174.150 3296.370 ;
        RECT 174.990 3295.720 179.210 3296.370 ;
        RECT 180.050 3295.720 184.270 3296.370 ;
        RECT 185.110 3295.720 189.330 3296.370 ;
        RECT 190.170 3295.720 194.390 3296.370 ;
        RECT 195.230 3295.720 199.450 3296.370 ;
        RECT 200.290 3295.720 204.510 3296.370 ;
        RECT 205.350 3295.720 209.570 3296.370 ;
        RECT 210.410 3295.720 214.630 3296.370 ;
        RECT 215.470 3295.720 219.690 3296.370 ;
        RECT 220.530 3295.720 224.750 3296.370 ;
        RECT 225.590 3295.720 229.810 3296.370 ;
        RECT 230.650 3295.720 234.870 3296.370 ;
        RECT 235.710 3295.720 239.930 3296.370 ;
        RECT 240.770 3295.720 244.990 3296.370 ;
        RECT 245.830 3295.720 250.050 3296.370 ;
        RECT 250.890 3295.720 255.110 3296.370 ;
        RECT 255.950 3295.720 260.170 3296.370 ;
        RECT 261.010 3295.720 265.230 3296.370 ;
        RECT 266.070 3295.720 270.290 3296.370 ;
        RECT 271.130 3295.720 275.350 3296.370 ;
        RECT 276.190 3295.720 280.410 3296.370 ;
        RECT 281.250 3295.720 285.470 3296.370 ;
        RECT 286.310 3295.720 290.530 3296.370 ;
        RECT 291.370 3295.720 295.590 3296.370 ;
        RECT 296.430 3295.720 300.650 3296.370 ;
        RECT 301.490 3295.720 305.710 3296.370 ;
        RECT 306.550 3295.720 310.770 3296.370 ;
        RECT 311.610 3295.720 315.830 3296.370 ;
        RECT 316.670 3295.720 320.890 3296.370 ;
        RECT 321.730 3295.720 325.950 3296.370 ;
        RECT 326.790 3295.720 331.010 3296.370 ;
        RECT 331.850 3295.720 336.070 3296.370 ;
        RECT 336.910 3295.720 341.130 3296.370 ;
        RECT 341.970 3295.720 346.190 3296.370 ;
        RECT 347.030 3295.720 351.250 3296.370 ;
        RECT 352.090 3295.720 356.310 3296.370 ;
        RECT 357.150 3295.720 361.370 3296.370 ;
        RECT 362.210 3295.720 366.430 3296.370 ;
        RECT 367.270 3295.720 371.490 3296.370 ;
        RECT 372.330 3295.720 376.550 3296.370 ;
        RECT 377.390 3295.720 381.610 3296.370 ;
        RECT 382.450 3295.720 386.670 3296.370 ;
        RECT 387.510 3295.720 391.730 3296.370 ;
        RECT 392.570 3295.720 396.790 3296.370 ;
        RECT 397.630 3295.720 401.850 3296.370 ;
        RECT 402.690 3295.720 406.910 3296.370 ;
        RECT 407.750 3295.720 411.970 3296.370 ;
        RECT 412.810 3295.720 417.030 3296.370 ;
        RECT 417.870 3295.720 422.090 3296.370 ;
        RECT 422.930 3295.720 427.150 3296.370 ;
        RECT 427.990 3295.720 432.210 3296.370 ;
        RECT 433.050 3295.720 437.270 3296.370 ;
        RECT 438.110 3295.720 442.330 3296.370 ;
        RECT 443.170 3295.720 447.390 3296.370 ;
        RECT 448.230 3295.720 452.450 3296.370 ;
        RECT 453.290 3295.720 457.510 3296.370 ;
        RECT 458.350 3295.720 462.570 3296.370 ;
        RECT 463.410 3295.720 467.630 3296.370 ;
        RECT 468.470 3295.720 472.690 3296.370 ;
        RECT 473.530 3295.720 477.750 3296.370 ;
        RECT 478.590 3295.720 482.810 3296.370 ;
        RECT 483.650 3295.720 487.870 3296.370 ;
        RECT 488.710 3295.720 492.930 3296.370 ;
        RECT 493.770 3295.720 497.990 3296.370 ;
        RECT 498.830 3295.720 503.050 3296.370 ;
        RECT 503.890 3295.720 508.110 3296.370 ;
        RECT 508.950 3295.720 513.170 3296.370 ;
        RECT 514.010 3295.720 518.230 3296.370 ;
        RECT 519.070 3295.720 523.290 3296.370 ;
        RECT 524.130 3295.720 528.350 3296.370 ;
        RECT 529.190 3295.720 533.410 3296.370 ;
        RECT 534.250 3295.720 538.470 3296.370 ;
        RECT 539.310 3295.720 543.530 3296.370 ;
        RECT 544.370 3295.720 548.590 3296.370 ;
        RECT 549.430 3295.720 553.650 3296.370 ;
        RECT 554.490 3295.720 558.710 3296.370 ;
        RECT 559.550 3295.720 563.770 3296.370 ;
        RECT 564.610 3295.720 568.830 3296.370 ;
        RECT 569.670 3295.720 573.890 3296.370 ;
        RECT 574.730 3295.720 578.950 3296.370 ;
        RECT 579.790 3295.720 584.010 3296.370 ;
        RECT 584.850 3295.720 589.070 3296.370 ;
        RECT 589.910 3295.720 594.130 3296.370 ;
        RECT 594.970 3295.720 599.190 3296.370 ;
        RECT 600.030 3295.720 604.250 3296.370 ;
        RECT 605.090 3295.720 609.310 3296.370 ;
        RECT 610.150 3295.720 614.370 3296.370 ;
        RECT 615.210 3295.720 619.430 3296.370 ;
        RECT 620.270 3295.720 624.490 3296.370 ;
        RECT 625.330 3295.720 629.550 3296.370 ;
        RECT 630.390 3295.720 634.610 3296.370 ;
        RECT 635.450 3295.720 639.670 3296.370 ;
        RECT 640.510 3295.720 644.730 3296.370 ;
        RECT 645.570 3295.720 649.790 3296.370 ;
        RECT 650.630 3295.720 654.850 3296.370 ;
        RECT 655.690 3295.720 659.910 3296.370 ;
        RECT 660.750 3295.720 664.970 3296.370 ;
        RECT 665.810 3295.720 670.030 3296.370 ;
        RECT 670.870 3295.720 675.090 3296.370 ;
        RECT 675.930 3295.720 680.150 3296.370 ;
        RECT 680.990 3295.720 685.210 3296.370 ;
        RECT 686.050 3295.720 690.270 3296.370 ;
        RECT 691.110 3295.720 695.330 3296.370 ;
        RECT 696.170 3295.720 700.390 3296.370 ;
        RECT 701.230 3295.720 705.450 3296.370 ;
        RECT 706.290 3295.720 710.510 3296.370 ;
        RECT 711.350 3295.720 715.570 3296.370 ;
        RECT 716.410 3295.720 720.630 3296.370 ;
        RECT 721.470 3295.720 725.690 3296.370 ;
        RECT 726.530 3295.720 730.750 3296.370 ;
        RECT 731.590 3295.720 735.810 3296.370 ;
        RECT 736.650 3295.720 740.870 3296.370 ;
        RECT 741.710 3295.720 745.930 3296.370 ;
        RECT 746.770 3295.720 750.990 3296.370 ;
        RECT 751.830 3295.720 756.050 3296.370 ;
        RECT 756.890 3295.720 761.110 3296.370 ;
        RECT 761.950 3295.720 766.170 3296.370 ;
        RECT 767.010 3295.720 771.230 3296.370 ;
        RECT 772.070 3295.720 776.290 3296.370 ;
        RECT 777.130 3295.720 781.350 3296.370 ;
        RECT 782.190 3295.720 786.410 3296.370 ;
        RECT 787.250 3295.720 791.470 3296.370 ;
        RECT 792.310 3295.720 796.530 3296.370 ;
        RECT 797.370 3295.720 801.590 3296.370 ;
        RECT 802.430 3295.720 806.650 3296.370 ;
        RECT 807.490 3295.720 811.710 3296.370 ;
        RECT 812.550 3295.720 816.770 3296.370 ;
        RECT 817.610 3295.720 821.830 3296.370 ;
        RECT 822.670 3295.720 826.890 3296.370 ;
        RECT 827.730 3295.720 831.950 3296.370 ;
        RECT 832.790 3295.720 837.010 3296.370 ;
        RECT 837.850 3295.720 842.070 3296.370 ;
        RECT 842.910 3295.720 847.130 3296.370 ;
        RECT 847.970 3295.720 852.190 3296.370 ;
        RECT 853.030 3295.720 857.250 3296.370 ;
        RECT 858.090 3295.720 862.310 3296.370 ;
        RECT 863.150 3295.720 867.370 3296.370 ;
        RECT 868.210 3295.720 872.430 3296.370 ;
        RECT 873.270 3295.720 877.490 3296.370 ;
        RECT 878.330 3295.720 882.550 3296.370 ;
        RECT 883.390 3295.720 887.610 3296.370 ;
        RECT 888.450 3295.720 892.670 3296.370 ;
        RECT 893.510 3295.720 897.730 3296.370 ;
        RECT 898.570 3295.720 902.790 3296.370 ;
        RECT 903.630 3295.720 907.850 3296.370 ;
        RECT 908.690 3295.720 912.910 3296.370 ;
        RECT 913.750 3295.720 917.970 3296.370 ;
        RECT 918.810 3295.720 923.030 3296.370 ;
        RECT 923.870 3295.720 928.090 3296.370 ;
        RECT 928.930 3295.720 933.150 3296.370 ;
        RECT 933.990 3295.720 938.210 3296.370 ;
        RECT 939.050 3295.720 943.270 3296.370 ;
        RECT 944.110 3295.720 948.330 3296.370 ;
        RECT 949.170 3295.720 953.390 3296.370 ;
        RECT 954.230 3295.720 958.450 3296.370 ;
        RECT 959.290 3295.720 963.510 3296.370 ;
        RECT 964.350 3295.720 968.570 3296.370 ;
        RECT 969.410 3295.720 973.630 3296.370 ;
        RECT 974.470 3295.720 978.690 3296.370 ;
        RECT 979.530 3295.720 983.750 3296.370 ;
        RECT 984.590 3295.720 988.810 3296.370 ;
        RECT 989.650 3295.720 993.870 3296.370 ;
        RECT 994.710 3295.720 998.930 3296.370 ;
        RECT 999.770 3295.720 1003.990 3296.370 ;
        RECT 1004.830 3295.720 1009.050 3296.370 ;
        RECT 1009.890 3295.720 1014.110 3296.370 ;
        RECT 1014.950 3295.720 1019.170 3296.370 ;
        RECT 1020.010 3295.720 1024.230 3296.370 ;
        RECT 1025.070 3295.720 1029.290 3296.370 ;
        RECT 1030.130 3295.720 1034.350 3296.370 ;
        RECT 1035.190 3295.720 1039.410 3296.370 ;
        RECT 1040.250 3295.720 1044.470 3296.370 ;
        RECT 1045.310 3295.720 1049.530 3296.370 ;
        RECT 1050.370 3295.720 1054.590 3296.370 ;
        RECT 1055.430 3295.720 1059.650 3296.370 ;
        RECT 1060.490 3295.720 1064.710 3296.370 ;
        RECT 1065.550 3295.720 1069.770 3296.370 ;
        RECT 1070.610 3295.720 1074.830 3296.370 ;
        RECT 1075.670 3295.720 1079.890 3296.370 ;
        RECT 1080.730 3295.720 1084.950 3296.370 ;
        RECT 1085.790 3295.720 1090.010 3296.370 ;
        RECT 1090.850 3295.720 1095.070 3296.370 ;
        RECT 1095.910 3295.720 1100.130 3296.370 ;
        RECT 1100.970 3295.720 1105.190 3296.370 ;
        RECT 1106.030 3295.720 1110.250 3296.370 ;
        RECT 1111.090 3295.720 1115.310 3296.370 ;
        RECT 1116.150 3295.720 1120.370 3296.370 ;
        RECT 1121.210 3295.720 1125.430 3296.370 ;
        RECT 1126.270 3295.720 1130.490 3296.370 ;
        RECT 1131.330 3295.720 1135.550 3296.370 ;
        RECT 1136.390 3295.720 1140.610 3296.370 ;
        RECT 1141.450 3295.720 1145.670 3296.370 ;
        RECT 1146.510 3295.720 1150.730 3296.370 ;
        RECT 1151.570 3295.720 1155.790 3296.370 ;
        RECT 1156.630 3295.720 1160.850 3296.370 ;
        RECT 1161.690 3295.720 1165.910 3296.370 ;
        RECT 1166.750 3295.720 1170.970 3296.370 ;
        RECT 1171.810 3295.720 1176.030 3296.370 ;
        RECT 1176.870 3295.720 1181.090 3296.370 ;
        RECT 1181.930 3295.720 1186.150 3296.370 ;
        RECT 1186.990 3295.720 1191.210 3296.370 ;
        RECT 1192.050 3295.720 1196.270 3296.370 ;
        RECT 1197.110 3295.720 1201.330 3296.370 ;
        RECT 1202.170 3295.720 1206.390 3296.370 ;
        RECT 1207.230 3295.720 1211.450 3296.370 ;
        RECT 1212.290 3295.720 1216.510 3296.370 ;
        RECT 1217.350 3295.720 1221.570 3296.370 ;
        RECT 1222.410 3295.720 1226.630 3296.370 ;
        RECT 1227.470 3295.720 1231.690 3296.370 ;
        RECT 1232.530 3295.720 1236.750 3296.370 ;
        RECT 1237.590 3295.720 1241.810 3296.370 ;
        RECT 1242.650 3295.720 1246.870 3296.370 ;
        RECT 1247.710 3295.720 1251.930 3296.370 ;
        RECT 1252.770 3295.720 1256.990 3296.370 ;
        RECT 1257.830 3295.720 1262.050 3296.370 ;
        RECT 1262.890 3295.720 1267.110 3296.370 ;
        RECT 1267.950 3295.720 1272.170 3296.370 ;
        RECT 1273.010 3295.720 1277.230 3296.370 ;
        RECT 1278.070 3295.720 1282.290 3296.370 ;
        RECT 1283.130 3295.720 1287.350 3296.370 ;
        RECT 1288.190 3295.720 1292.410 3296.370 ;
        RECT 1293.250 3295.720 1297.470 3296.370 ;
        RECT 1298.310 3295.720 1302.530 3296.370 ;
        RECT 1303.370 3295.720 1307.590 3296.370 ;
        RECT 1308.430 3295.720 1312.650 3296.370 ;
        RECT 1313.490 3295.720 1317.710 3296.370 ;
        RECT 1318.550 3295.720 1322.770 3296.370 ;
        RECT 1323.610 3295.720 1327.830 3296.370 ;
        RECT 1328.670 3295.720 1332.890 3296.370 ;
        RECT 1333.730 3295.720 1337.950 3296.370 ;
        RECT 1338.790 3295.720 1343.010 3296.370 ;
        RECT 1343.850 3295.720 1348.070 3296.370 ;
        RECT 1348.910 3295.720 1353.130 3296.370 ;
        RECT 1353.970 3295.720 1358.190 3296.370 ;
        RECT 1359.030 3295.720 1363.250 3296.370 ;
        RECT 1364.090 3295.720 1368.310 3296.370 ;
        RECT 1369.150 3295.720 1373.370 3296.370 ;
        RECT 1374.210 3295.720 1378.430 3296.370 ;
        RECT 1379.270 3295.720 1383.490 3296.370 ;
        RECT 1384.330 3295.720 1388.550 3296.370 ;
        RECT 1389.390 3295.720 1393.610 3296.370 ;
        RECT 1394.450 3295.720 1398.670 3296.370 ;
        RECT 1399.510 3295.720 1403.730 3296.370 ;
        RECT 1404.570 3295.720 1408.790 3296.370 ;
        RECT 1409.630 3295.720 1413.850 3296.370 ;
        RECT 1414.690 3295.720 1418.910 3296.370 ;
        RECT 1419.750 3295.720 1423.970 3296.370 ;
        RECT 1424.810 3295.720 1429.030 3296.370 ;
        RECT 1429.870 3295.720 1434.090 3296.370 ;
        RECT 1434.930 3295.720 1439.150 3296.370 ;
        RECT 1439.990 3295.720 1444.210 3296.370 ;
        RECT 1445.050 3295.720 1449.270 3296.370 ;
        RECT 1450.110 3295.720 1454.330 3296.370 ;
        RECT 1455.170 3295.720 1459.390 3296.370 ;
        RECT 1460.230 3295.720 1464.450 3296.370 ;
        RECT 1465.290 3295.720 1469.510 3296.370 ;
        RECT 1470.350 3295.720 1474.570 3296.370 ;
        RECT 1475.410 3295.720 1479.630 3296.370 ;
        RECT 1480.470 3295.720 1484.690 3296.370 ;
        RECT 1485.530 3295.720 1489.750 3296.370 ;
        RECT 1490.590 3295.720 1494.810 3296.370 ;
        RECT 1495.650 3295.720 1499.870 3296.370 ;
        RECT 1500.710 3295.720 1504.930 3296.370 ;
        RECT 1505.770 3295.720 1509.990 3296.370 ;
        RECT 1510.830 3295.720 1515.050 3296.370 ;
        RECT 1515.890 3295.720 1520.110 3296.370 ;
        RECT 1520.950 3295.720 1525.170 3296.370 ;
        RECT 1526.010 3295.720 1530.230 3296.370 ;
        RECT 1531.070 3295.720 1535.290 3296.370 ;
        RECT 1536.130 3295.720 1540.350 3296.370 ;
        RECT 1541.190 3295.720 1545.410 3296.370 ;
        RECT 1546.250 3295.720 1550.470 3296.370 ;
        RECT 1551.310 3295.720 1555.530 3296.370 ;
        RECT 1556.370 3295.720 1560.590 3296.370 ;
        RECT 1561.430 3295.720 1565.650 3296.370 ;
        RECT 1566.490 3295.720 1570.710 3296.370 ;
        RECT 1571.550 3295.720 1575.770 3296.370 ;
        RECT 1576.610 3295.720 1580.830 3296.370 ;
        RECT 1581.670 3295.720 1585.890 3296.370 ;
        RECT 1586.730 3295.720 1590.950 3296.370 ;
        RECT 1591.790 3295.720 1596.010 3296.370 ;
        RECT 1596.850 3295.720 1601.070 3296.370 ;
        RECT 1601.910 3295.720 1606.130 3296.370 ;
        RECT 1606.970 3295.720 1611.190 3296.370 ;
        RECT 1612.030 3295.720 1616.250 3296.370 ;
        RECT 1617.090 3295.720 1621.310 3296.370 ;
        RECT 1622.150 3295.720 1626.370 3296.370 ;
        RECT 1627.210 3295.720 1631.430 3296.370 ;
        RECT 1632.270 3295.720 1636.490 3296.370 ;
        RECT 1637.330 3295.720 1641.550 3296.370 ;
        RECT 1642.390 3295.720 1646.610 3296.370 ;
        RECT 1647.450 3295.720 1651.670 3296.370 ;
        RECT 1652.510 3295.720 1656.730 3296.370 ;
        RECT 1657.570 3295.720 1661.790 3296.370 ;
        RECT 1662.630 3295.720 1666.850 3296.370 ;
        RECT 1667.690 3295.720 1671.910 3296.370 ;
        RECT 1672.750 3295.720 1676.970 3296.370 ;
        RECT 1677.810 3295.720 1682.030 3296.370 ;
        RECT 1682.870 3295.720 1687.090 3296.370 ;
        RECT 1687.930 3295.720 1692.150 3296.370 ;
        RECT 1692.990 3295.720 1697.210 3296.370 ;
        RECT 1698.050 3295.720 1702.270 3296.370 ;
        RECT 1703.110 3295.720 1707.330 3296.370 ;
        RECT 1708.170 3295.720 1712.390 3296.370 ;
        RECT 1713.230 3295.720 1717.450 3296.370 ;
        RECT 1718.290 3295.720 1722.510 3296.370 ;
        RECT 1723.350 3295.720 1727.570 3296.370 ;
        RECT 1728.410 3295.720 1732.630 3296.370 ;
        RECT 1733.470 3295.720 1737.690 3296.370 ;
        RECT 1738.530 3295.720 1742.750 3296.370 ;
        RECT 1743.590 3295.720 1747.810 3296.370 ;
        RECT 1748.650 3295.720 1752.870 3296.370 ;
        RECT 1753.710 3295.720 1757.930 3296.370 ;
        RECT 1758.770 3295.720 1762.990 3296.370 ;
        RECT 1763.830 3295.720 1768.050 3296.370 ;
        RECT 1768.890 3295.720 1773.110 3296.370 ;
        RECT 1773.950 3295.720 1778.170 3296.370 ;
        RECT 1779.010 3295.720 1783.230 3296.370 ;
        RECT 1784.070 3295.720 1788.290 3296.370 ;
        RECT 1789.130 3295.720 1793.350 3296.370 ;
        RECT 1794.190 3295.720 1798.410 3296.370 ;
        RECT 1799.250 3295.720 1803.470 3296.370 ;
        RECT 1804.310 3295.720 1808.530 3296.370 ;
        RECT 1809.370 3295.720 1813.590 3296.370 ;
        RECT 1814.430 3295.720 1818.650 3296.370 ;
        RECT 1819.490 3295.720 1823.710 3296.370 ;
        RECT 1824.550 3295.720 1828.770 3296.370 ;
        RECT 1829.610 3295.720 1833.830 3296.370 ;
        RECT 1834.670 3295.720 1838.890 3296.370 ;
        RECT 1839.730 3295.720 1843.950 3296.370 ;
        RECT 1844.790 3295.720 1849.010 3296.370 ;
        RECT 1849.850 3295.720 1854.070 3296.370 ;
        RECT 1854.910 3295.720 1859.130 3296.370 ;
        RECT 1859.970 3295.720 1864.190 3296.370 ;
        RECT 1865.030 3295.720 1869.250 3296.370 ;
        RECT 1870.090 3295.720 1874.310 3296.370 ;
        RECT 1875.150 3295.720 1879.370 3296.370 ;
        RECT 1880.210 3295.720 1884.430 3296.370 ;
        RECT 1885.270 3295.720 1889.490 3296.370 ;
        RECT 1890.330 3295.720 1894.550 3296.370 ;
        RECT 1895.390 3295.720 1899.610 3296.370 ;
        RECT 1900.450 3295.720 1904.670 3296.370 ;
        RECT 1905.510 3295.720 1909.730 3296.370 ;
        RECT 1910.570 3295.720 1914.790 3296.370 ;
        RECT 1915.630 3295.720 1919.850 3296.370 ;
        RECT 1920.690 3295.720 1924.910 3296.370 ;
        RECT 1925.750 3295.720 1929.970 3296.370 ;
        RECT 1930.810 3295.720 1935.030 3296.370 ;
        RECT 1935.870 3295.720 1940.090 3296.370 ;
        RECT 1940.930 3295.720 1945.150 3296.370 ;
        RECT 1945.990 3295.720 1950.210 3296.370 ;
        RECT 1951.050 3295.720 1955.270 3296.370 ;
        RECT 1956.110 3295.720 1960.330 3296.370 ;
        RECT 1961.170 3295.720 1965.390 3296.370 ;
        RECT 1966.230 3295.720 1970.450 3296.370 ;
        RECT 1971.290 3295.720 1975.510 3296.370 ;
        RECT 1976.350 3295.720 1980.570 3296.370 ;
        RECT 1981.410 3295.720 1985.630 3296.370 ;
        RECT 1986.470 3295.720 1990.690 3296.370 ;
        RECT 1991.530 3295.720 1995.750 3296.370 ;
        RECT 1996.590 3295.720 2000.810 3296.370 ;
        RECT 2001.650 3295.720 2005.870 3296.370 ;
        RECT 2006.710 3295.720 2010.930 3296.370 ;
        RECT 2011.770 3295.720 2015.990 3296.370 ;
        RECT 2016.830 3295.720 2021.050 3296.370 ;
        RECT 2021.890 3295.720 2026.110 3296.370 ;
        RECT 2026.950 3295.720 2092.910 3296.370 ;
        RECT 4.690 4.280 2092.910 3295.720 ;
        RECT 4.690 4.000 10.850 4.280 ;
        RECT 11.690 4.000 30.630 4.280 ;
        RECT 31.470 4.000 50.410 4.280 ;
        RECT 51.250 4.000 70.190 4.280 ;
        RECT 71.030 4.000 89.970 4.280 ;
        RECT 90.810 4.000 109.750 4.280 ;
        RECT 110.590 4.000 129.530 4.280 ;
        RECT 130.370 4.000 149.310 4.280 ;
        RECT 150.150 4.000 169.090 4.280 ;
        RECT 169.930 4.000 188.870 4.280 ;
        RECT 189.710 4.000 208.650 4.280 ;
        RECT 209.490 4.000 228.430 4.280 ;
        RECT 229.270 4.000 248.210 4.280 ;
        RECT 249.050 4.000 267.990 4.280 ;
        RECT 268.830 4.000 287.770 4.280 ;
        RECT 288.610 4.000 307.550 4.280 ;
        RECT 308.390 4.000 327.330 4.280 ;
        RECT 328.170 4.000 347.110 4.280 ;
        RECT 347.950 4.000 366.890 4.280 ;
        RECT 367.730 4.000 386.670 4.280 ;
        RECT 387.510 4.000 406.450 4.280 ;
        RECT 407.290 4.000 426.230 4.280 ;
        RECT 427.070 4.000 446.010 4.280 ;
        RECT 446.850 4.000 465.790 4.280 ;
        RECT 466.630 4.000 485.570 4.280 ;
        RECT 486.410 4.000 505.350 4.280 ;
        RECT 506.190 4.000 525.130 4.280 ;
        RECT 525.970 4.000 544.910 4.280 ;
        RECT 545.750 4.000 564.690 4.280 ;
        RECT 565.530 4.000 584.470 4.280 ;
        RECT 585.310 4.000 604.250 4.280 ;
        RECT 605.090 4.000 624.030 4.280 ;
        RECT 624.870 4.000 643.810 4.280 ;
        RECT 644.650 4.000 663.590 4.280 ;
        RECT 664.430 4.000 683.370 4.280 ;
        RECT 684.210 4.000 703.150 4.280 ;
        RECT 703.990 4.000 722.930 4.280 ;
        RECT 723.770 4.000 742.710 4.280 ;
        RECT 743.550 4.000 762.490 4.280 ;
        RECT 763.330 4.000 782.270 4.280 ;
        RECT 783.110 4.000 802.050 4.280 ;
        RECT 802.890 4.000 821.830 4.280 ;
        RECT 822.670 4.000 841.610 4.280 ;
        RECT 842.450 4.000 861.390 4.280 ;
        RECT 862.230 4.000 881.170 4.280 ;
        RECT 882.010 4.000 900.950 4.280 ;
        RECT 901.790 4.000 920.730 4.280 ;
        RECT 921.570 4.000 940.510 4.280 ;
        RECT 941.350 4.000 960.290 4.280 ;
        RECT 961.130 4.000 980.070 4.280 ;
        RECT 980.910 4.000 999.850 4.280 ;
        RECT 1000.690 4.000 1019.630 4.280 ;
        RECT 1020.470 4.000 1039.410 4.280 ;
        RECT 1040.250 4.000 1059.190 4.280 ;
        RECT 1060.030 4.000 1078.970 4.280 ;
        RECT 1079.810 4.000 1098.750 4.280 ;
        RECT 1099.590 4.000 1118.530 4.280 ;
        RECT 1119.370 4.000 1138.310 4.280 ;
        RECT 1139.150 4.000 1158.090 4.280 ;
        RECT 1158.930 4.000 1177.870 4.280 ;
        RECT 1178.710 4.000 1197.650 4.280 ;
        RECT 1198.490 4.000 1217.430 4.280 ;
        RECT 1218.270 4.000 1237.210 4.280 ;
        RECT 1238.050 4.000 1256.990 4.280 ;
        RECT 1257.830 4.000 1276.770 4.280 ;
        RECT 1277.610 4.000 1296.550 4.280 ;
        RECT 1297.390 4.000 1316.330 4.280 ;
        RECT 1317.170 4.000 1336.110 4.280 ;
        RECT 1336.950 4.000 1355.890 4.280 ;
        RECT 1356.730 4.000 1375.670 4.280 ;
        RECT 1376.510 4.000 1395.450 4.280 ;
        RECT 1396.290 4.000 1415.230 4.280 ;
        RECT 1416.070 4.000 1435.010 4.280 ;
        RECT 1435.850 4.000 1454.790 4.280 ;
        RECT 1455.630 4.000 1474.570 4.280 ;
        RECT 1475.410 4.000 1494.350 4.280 ;
        RECT 1495.190 4.000 1514.130 4.280 ;
        RECT 1514.970 4.000 1533.910 4.280 ;
        RECT 1534.750 4.000 1553.690 4.280 ;
        RECT 1554.530 4.000 1573.470 4.280 ;
        RECT 1574.310 4.000 1593.250 4.280 ;
        RECT 1594.090 4.000 1613.030 4.280 ;
        RECT 1613.870 4.000 1632.810 4.280 ;
        RECT 1633.650 4.000 1652.590 4.280 ;
        RECT 1653.430 4.000 1672.370 4.280 ;
        RECT 1673.210 4.000 1692.150 4.280 ;
        RECT 1692.990 4.000 1711.930 4.280 ;
        RECT 1712.770 4.000 1731.710 4.280 ;
        RECT 1732.550 4.000 1751.490 4.280 ;
        RECT 1752.330 4.000 1771.270 4.280 ;
        RECT 1772.110 4.000 1791.050 4.280 ;
        RECT 1791.890 4.000 1810.830 4.280 ;
        RECT 1811.670 4.000 1830.610 4.280 ;
        RECT 1831.450 4.000 1850.390 4.280 ;
        RECT 1851.230 4.000 1870.170 4.280 ;
        RECT 1871.010 4.000 1889.950 4.280 ;
        RECT 1890.790 4.000 1909.730 4.280 ;
        RECT 1910.570 4.000 1929.510 4.280 ;
        RECT 1930.350 4.000 1949.290 4.280 ;
        RECT 1950.130 4.000 1969.070 4.280 ;
        RECT 1969.910 4.000 1988.850 4.280 ;
        RECT 1989.690 4.000 2008.630 4.280 ;
        RECT 2009.470 4.000 2028.410 4.280 ;
        RECT 2029.250 4.000 2048.190 4.280 ;
        RECT 2049.030 4.000 2067.970 4.280 ;
        RECT 2068.810 4.000 2087.750 4.280 ;
        RECT 2088.590 4.000 2092.910 4.280 ;
      LAYER met3 ;
        RECT 4.000 3229.680 2096.000 3288.645 ;
        RECT 4.400 3228.280 2095.600 3229.680 ;
        RECT 4.000 3092.320 2096.000 3228.280 ;
        RECT 4.400 3090.920 2095.600 3092.320 ;
        RECT 4.000 2954.960 2096.000 3090.920 ;
        RECT 4.400 2953.560 2095.600 2954.960 ;
        RECT 4.000 2817.600 2096.000 2953.560 ;
        RECT 4.400 2816.200 2095.600 2817.600 ;
        RECT 4.000 2680.240 2096.000 2816.200 ;
        RECT 4.400 2678.840 2095.600 2680.240 ;
        RECT 4.000 2542.880 2096.000 2678.840 ;
        RECT 4.400 2541.480 2095.600 2542.880 ;
        RECT 4.000 2405.520 2096.000 2541.480 ;
        RECT 4.400 2404.120 2095.600 2405.520 ;
        RECT 4.000 2268.160 2096.000 2404.120 ;
        RECT 4.400 2266.760 2095.600 2268.160 ;
        RECT 4.000 2130.800 2096.000 2266.760 ;
        RECT 4.400 2129.400 2095.600 2130.800 ;
        RECT 4.000 1993.440 2096.000 2129.400 ;
        RECT 4.400 1992.040 2095.600 1993.440 ;
        RECT 4.000 1856.080 2096.000 1992.040 ;
        RECT 4.400 1854.680 2095.600 1856.080 ;
        RECT 4.000 1718.720 2096.000 1854.680 ;
        RECT 4.400 1717.320 2095.600 1718.720 ;
        RECT 4.000 1581.360 2096.000 1717.320 ;
        RECT 4.400 1579.960 2095.600 1581.360 ;
        RECT 4.000 1444.000 2096.000 1579.960 ;
        RECT 4.400 1442.600 2095.600 1444.000 ;
        RECT 4.000 1306.640 2096.000 1442.600 ;
        RECT 4.400 1305.240 2095.600 1306.640 ;
        RECT 4.000 1169.280 2096.000 1305.240 ;
        RECT 4.400 1167.880 2095.600 1169.280 ;
        RECT 4.000 1031.920 2096.000 1167.880 ;
        RECT 4.400 1030.520 2095.600 1031.920 ;
        RECT 4.000 894.560 2096.000 1030.520 ;
        RECT 4.400 893.160 2095.600 894.560 ;
        RECT 4.000 757.200 2096.000 893.160 ;
        RECT 4.400 755.800 2095.600 757.200 ;
        RECT 4.000 619.840 2096.000 755.800 ;
        RECT 4.400 618.440 2095.600 619.840 ;
        RECT 4.000 482.480 2096.000 618.440 ;
        RECT 4.400 481.080 2095.600 482.480 ;
        RECT 4.000 345.120 2096.000 481.080 ;
        RECT 4.400 343.720 2095.600 345.120 ;
        RECT 4.000 207.760 2096.000 343.720 ;
        RECT 4.400 206.360 2095.600 207.760 ;
        RECT 4.000 70.400 2096.000 206.360 ;
        RECT 4.400 69.000 2095.600 70.400 ;
        RECT 4.000 10.715 2096.000 69.000 ;
      LAYER met4 ;
        RECT 187.975 191.935 251.320 3286.945 ;
        RECT 253.720 191.935 254.620 3286.945 ;
        RECT 257.020 191.935 321.320 3286.945 ;
        RECT 323.720 191.935 324.620 3286.945 ;
        RECT 327.020 191.935 391.320 3286.945 ;
        RECT 393.720 191.935 394.620 3286.945 ;
        RECT 397.020 3087.180 461.320 3286.945 ;
        RECT 463.720 3087.180 464.620 3286.945 ;
        RECT 397.020 3010.740 464.620 3087.180 ;
        RECT 397.020 2889.785 461.320 3010.740 ;
        RECT 463.720 2889.785 464.620 3010.740 ;
        RECT 467.020 2889.785 531.320 3286.945 ;
        RECT 397.020 2836.695 531.320 2889.785 ;
        RECT 397.020 2810.740 464.620 2836.695 ;
        RECT 397.020 2287.180 461.320 2810.740 ;
        RECT 463.720 2698.060 464.620 2810.740 ;
        RECT 467.020 2698.060 531.320 2836.695 ;
        RECT 463.720 2610.740 531.320 2698.060 ;
        RECT 463.720 2287.180 464.620 2610.740 ;
        RECT 397.020 2210.740 464.620 2287.180 ;
        RECT 397.020 1687.180 461.320 2210.740 ;
        RECT 463.720 2098.060 464.620 2210.740 ;
        RECT 467.020 2098.060 531.320 2610.740 ;
        RECT 463.720 2010.740 531.320 2098.060 ;
        RECT 463.720 1687.180 464.620 2010.740 ;
        RECT 397.020 1610.740 464.620 1687.180 ;
        RECT 397.020 1087.180 461.320 1610.740 ;
        RECT 463.720 1498.060 464.620 1610.740 ;
        RECT 467.020 1498.060 531.320 2010.740 ;
        RECT 463.720 1410.740 531.320 1498.060 ;
        RECT 463.720 1087.180 464.620 1410.740 ;
        RECT 397.020 1010.740 464.620 1087.180 ;
        RECT 397.020 487.180 461.320 1010.740 ;
        RECT 463.720 898.060 464.620 1010.740 ;
        RECT 467.020 898.060 531.320 1410.740 ;
        RECT 463.720 810.740 531.320 898.060 ;
        RECT 463.720 487.180 464.620 810.740 ;
        RECT 397.020 410.740 464.620 487.180 ;
        RECT 397.020 287.180 461.320 410.740 ;
        RECT 463.720 287.180 464.620 410.740 ;
        RECT 397.020 210.740 464.620 287.180 ;
        RECT 397.020 191.935 461.320 210.740 ;
        RECT 463.720 191.935 464.620 210.740 ;
        RECT 467.020 191.935 531.320 810.740 ;
        RECT 533.720 191.935 534.620 3286.945 ;
        RECT 537.020 191.935 601.320 3286.945 ;
        RECT 603.720 2683.665 604.620 3286.945 ;
        RECT 607.020 2887.180 671.320 3286.945 ;
        RECT 673.720 2887.180 674.620 3286.945 ;
        RECT 607.020 2880.265 674.620 2887.180 ;
        RECT 677.020 2880.265 741.320 3286.945 ;
        RECT 607.020 2812.895 741.320 2880.265 ;
        RECT 607.020 2810.740 674.620 2812.895 ;
        RECT 607.020 2687.180 671.320 2810.740 ;
        RECT 673.720 2687.180 674.620 2810.740 ;
        RECT 607.020 2683.665 674.620 2687.180 ;
        RECT 677.020 2683.665 741.320 2812.895 ;
        RECT 603.720 2612.215 741.320 2683.665 ;
        RECT 603.720 2283.665 604.620 2612.215 ;
        RECT 607.020 2610.740 674.620 2612.215 ;
        RECT 607.020 2287.180 671.320 2610.740 ;
        RECT 673.720 2287.180 674.620 2610.740 ;
        RECT 607.020 2283.665 674.620 2287.180 ;
        RECT 677.020 2283.665 741.320 2612.215 ;
        RECT 603.720 2206.095 741.320 2283.665 ;
        RECT 603.720 2083.665 604.620 2206.095 ;
        RECT 607.020 2087.180 671.320 2206.095 ;
        RECT 673.720 2087.180 674.620 2206.095 ;
        RECT 607.020 2083.665 674.620 2087.180 ;
        RECT 677.020 2083.665 741.320 2206.095 ;
        RECT 603.720 2012.215 741.320 2083.665 ;
        RECT 603.720 1683.665 604.620 2012.215 ;
        RECT 607.020 2010.740 674.620 2012.215 ;
        RECT 607.020 1687.180 671.320 2010.740 ;
        RECT 673.720 1687.180 674.620 2010.740 ;
        RECT 607.020 1683.665 674.620 1687.180 ;
        RECT 677.020 1683.665 741.320 2012.215 ;
        RECT 603.720 1606.095 741.320 1683.665 ;
        RECT 603.720 1483.665 604.620 1606.095 ;
        RECT 607.020 1487.180 671.320 1606.095 ;
        RECT 673.720 1487.180 674.620 1606.095 ;
        RECT 607.020 1483.665 674.620 1487.180 ;
        RECT 677.020 1483.665 741.320 1606.095 ;
        RECT 603.720 1412.215 741.320 1483.665 ;
        RECT 603.720 1083.665 604.620 1412.215 ;
        RECT 607.020 1410.740 674.620 1412.215 ;
        RECT 607.020 1087.180 671.320 1410.740 ;
        RECT 673.720 1087.180 674.620 1410.740 ;
        RECT 607.020 1083.665 674.620 1087.180 ;
        RECT 677.020 1083.665 741.320 1412.215 ;
        RECT 603.720 1006.095 741.320 1083.665 ;
        RECT 603.720 883.665 604.620 1006.095 ;
        RECT 607.020 887.180 671.320 1006.095 ;
        RECT 673.720 887.180 674.620 1006.095 ;
        RECT 607.020 883.665 674.620 887.180 ;
        RECT 677.020 883.665 741.320 1006.095 ;
        RECT 603.720 812.215 741.320 883.665 ;
        RECT 603.720 191.935 604.620 812.215 ;
        RECT 607.020 810.740 674.620 812.215 ;
        RECT 607.020 487.180 671.320 810.740 ;
        RECT 673.720 487.180 674.620 810.740 ;
        RECT 607.020 471.425 674.620 487.180 ;
        RECT 677.020 471.425 741.320 812.215 ;
        RECT 607.020 427.855 741.320 471.425 ;
        RECT 607.020 410.740 674.620 427.855 ;
        RECT 607.020 191.935 671.320 410.740 ;
        RECT 673.720 191.935 674.620 410.740 ;
        RECT 677.020 191.935 741.320 427.855 ;
        RECT 743.720 191.935 744.620 3286.945 ;
        RECT 747.020 2889.785 811.320 3286.945 ;
        RECT 813.720 3087.180 814.620 3286.945 ;
        RECT 817.020 3087.180 881.320 3286.945 ;
        RECT 883.720 3087.180 884.620 3286.945 ;
        RECT 813.720 3010.740 884.620 3087.180 ;
        RECT 813.720 2889.785 814.620 3010.740 ;
        RECT 817.020 2889.785 881.320 3010.740 ;
        RECT 883.720 2889.785 884.620 3010.740 ;
        RECT 887.020 2889.785 951.320 3286.945 ;
        RECT 747.020 2836.695 951.320 2889.785 ;
        RECT 747.020 191.935 811.320 2836.695 ;
        RECT 813.720 2810.740 884.620 2836.695 ;
        RECT 813.720 2698.060 814.620 2810.740 ;
        RECT 817.020 2698.060 881.320 2810.740 ;
        RECT 813.720 2687.065 881.320 2698.060 ;
        RECT 883.720 2687.065 884.620 2810.740 ;
        RECT 887.020 2687.065 951.320 2836.695 ;
        RECT 813.720 2616.975 951.320 2687.065 ;
        RECT 813.720 2610.740 881.320 2616.975 ;
        RECT 813.720 2287.180 814.620 2610.740 ;
        RECT 817.020 2287.180 881.320 2610.740 ;
        RECT 883.720 2287.180 884.620 2616.975 ;
        RECT 813.720 2210.740 884.620 2287.180 ;
        RECT 813.720 2098.060 814.620 2210.740 ;
        RECT 817.020 2098.060 881.320 2210.740 ;
        RECT 813.720 2087.065 881.320 2098.060 ;
        RECT 883.720 2087.065 884.620 2210.740 ;
        RECT 887.020 2087.065 951.320 2616.975 ;
        RECT 813.720 2016.975 951.320 2087.065 ;
        RECT 813.720 2010.740 881.320 2016.975 ;
        RECT 813.720 1687.180 814.620 2010.740 ;
        RECT 817.020 1687.180 881.320 2010.740 ;
        RECT 883.720 1687.180 884.620 2016.975 ;
        RECT 813.720 1610.740 884.620 1687.180 ;
        RECT 813.720 1498.060 814.620 1610.740 ;
        RECT 817.020 1498.060 881.320 1610.740 ;
        RECT 813.720 1487.065 881.320 1498.060 ;
        RECT 883.720 1487.065 884.620 1610.740 ;
        RECT 887.020 1487.065 951.320 2016.975 ;
        RECT 813.720 1416.975 951.320 1487.065 ;
        RECT 813.720 1410.740 881.320 1416.975 ;
        RECT 813.720 1087.180 814.620 1410.740 ;
        RECT 817.020 1087.180 881.320 1410.740 ;
        RECT 883.720 1087.180 884.620 1416.975 ;
        RECT 813.720 1010.740 884.620 1087.180 ;
        RECT 813.720 898.060 814.620 1010.740 ;
        RECT 817.020 898.060 881.320 1010.740 ;
        RECT 813.720 887.065 881.320 898.060 ;
        RECT 883.720 887.065 884.620 1010.740 ;
        RECT 887.020 887.065 951.320 1416.975 ;
        RECT 813.720 816.975 951.320 887.065 ;
        RECT 813.720 810.740 881.320 816.975 ;
        RECT 813.720 487.180 814.620 810.740 ;
        RECT 817.020 487.180 881.320 810.740 ;
        RECT 883.720 487.180 884.620 816.975 ;
        RECT 813.720 436.745 884.620 487.180 ;
        RECT 887.020 436.745 951.320 816.975 ;
        RECT 813.720 427.175 951.320 436.745 ;
        RECT 813.720 410.740 884.620 427.175 ;
        RECT 813.720 287.180 814.620 410.740 ;
        RECT 817.020 287.180 881.320 410.740 ;
        RECT 883.720 287.180 884.620 410.740 ;
        RECT 813.720 210.740 884.620 287.180 ;
        RECT 813.720 191.935 814.620 210.740 ;
        RECT 817.020 191.935 881.320 210.740 ;
        RECT 883.720 191.935 884.620 210.740 ;
        RECT 887.020 191.935 951.320 427.175 ;
        RECT 953.720 191.935 954.620 3286.945 ;
        RECT 957.020 2683.665 1021.320 3286.945 ;
        RECT 1023.720 2887.180 1024.620 3286.945 ;
        RECT 1027.020 2887.180 1091.320 3286.945 ;
        RECT 1093.720 2887.180 1094.620 3286.945 ;
        RECT 1097.020 2887.180 1161.320 3286.945 ;
        RECT 1023.720 2810.740 1161.320 2887.180 ;
        RECT 1023.720 2687.180 1024.620 2810.740 ;
        RECT 1027.020 2687.180 1091.320 2810.740 ;
        RECT 1093.720 2687.180 1094.620 2810.740 ;
        RECT 1097.020 2687.180 1161.320 2810.740 ;
        RECT 1023.720 2683.665 1161.320 2687.180 ;
        RECT 957.020 2612.215 1161.320 2683.665 ;
        RECT 957.020 2283.665 1021.320 2612.215 ;
        RECT 1023.720 2610.740 1161.320 2612.215 ;
        RECT 1023.720 2287.180 1024.620 2610.740 ;
        RECT 1027.020 2287.180 1091.320 2610.740 ;
        RECT 1093.720 2287.180 1094.620 2610.740 ;
        RECT 1097.020 2287.180 1161.320 2610.740 ;
        RECT 1023.720 2283.665 1161.320 2287.180 ;
        RECT 957.020 2206.095 1161.320 2283.665 ;
        RECT 957.020 2083.665 1021.320 2206.095 ;
        RECT 1023.720 2087.180 1024.620 2206.095 ;
        RECT 1027.020 2087.180 1091.320 2206.095 ;
        RECT 1093.720 2087.180 1094.620 2206.095 ;
        RECT 1097.020 2087.180 1161.320 2206.095 ;
        RECT 1023.720 2083.665 1161.320 2087.180 ;
        RECT 957.020 2012.215 1161.320 2083.665 ;
        RECT 957.020 1683.665 1021.320 2012.215 ;
        RECT 1023.720 2010.740 1161.320 2012.215 ;
        RECT 1023.720 1687.180 1024.620 2010.740 ;
        RECT 1027.020 1687.180 1091.320 2010.740 ;
        RECT 1093.720 1687.180 1094.620 2010.740 ;
        RECT 1097.020 1687.180 1161.320 2010.740 ;
        RECT 1023.720 1683.665 1161.320 1687.180 ;
        RECT 957.020 1606.095 1161.320 1683.665 ;
        RECT 957.020 1483.665 1021.320 1606.095 ;
        RECT 1023.720 1487.180 1024.620 1606.095 ;
        RECT 1027.020 1487.180 1091.320 1606.095 ;
        RECT 1093.720 1487.180 1094.620 1606.095 ;
        RECT 1097.020 1487.180 1161.320 1606.095 ;
        RECT 1023.720 1483.665 1161.320 1487.180 ;
        RECT 957.020 1412.215 1161.320 1483.665 ;
        RECT 957.020 1083.665 1021.320 1412.215 ;
        RECT 1023.720 1410.740 1161.320 1412.215 ;
        RECT 1023.720 1087.180 1024.620 1410.740 ;
        RECT 1027.020 1087.180 1091.320 1410.740 ;
        RECT 1093.720 1087.180 1094.620 1410.740 ;
        RECT 1097.020 1087.180 1161.320 1410.740 ;
        RECT 1023.720 1083.665 1161.320 1087.180 ;
        RECT 957.020 1006.095 1161.320 1083.665 ;
        RECT 957.020 883.665 1021.320 1006.095 ;
        RECT 1023.720 887.180 1024.620 1006.095 ;
        RECT 1027.020 887.180 1091.320 1006.095 ;
        RECT 1093.720 887.180 1094.620 1006.095 ;
        RECT 1097.020 887.180 1161.320 1006.095 ;
        RECT 1023.720 883.665 1161.320 887.180 ;
        RECT 957.020 812.215 1161.320 883.665 ;
        RECT 957.020 191.935 1021.320 812.215 ;
        RECT 1023.720 810.740 1161.320 812.215 ;
        RECT 1023.720 487.180 1024.620 810.740 ;
        RECT 1027.020 487.180 1091.320 810.740 ;
        RECT 1093.720 487.180 1094.620 810.740 ;
        RECT 1097.020 487.180 1161.320 810.740 ;
        RECT 1023.720 410.740 1161.320 487.180 ;
        RECT 1023.720 191.935 1024.620 410.740 ;
        RECT 1027.020 191.935 1091.320 410.740 ;
        RECT 1093.720 191.935 1094.620 410.740 ;
        RECT 1097.020 191.935 1161.320 410.740 ;
        RECT 1163.720 191.935 1164.620 3286.945 ;
        RECT 1167.020 2889.785 1231.320 3286.945 ;
        RECT 1233.720 2889.785 1234.620 3286.945 ;
        RECT 1237.020 2889.785 1301.320 3286.945 ;
        RECT 1167.020 2836.695 1301.320 2889.785 ;
        RECT 1167.020 2276.865 1231.320 2836.695 ;
        RECT 1233.720 2276.865 1234.620 2836.695 ;
        RECT 1237.020 2698.060 1301.320 2836.695 ;
        RECT 1303.720 2698.060 1304.620 3286.945 ;
        RECT 1307.020 2698.060 1371.320 3286.945 ;
        RECT 1237.020 2610.740 1371.320 2698.060 ;
        RECT 1237.020 2276.865 1301.320 2610.740 ;
        RECT 1167.020 2230.575 1301.320 2276.865 ;
        RECT 1167.020 1676.865 1231.320 2230.575 ;
        RECT 1233.720 1676.865 1234.620 2230.575 ;
        RECT 1237.020 2098.060 1301.320 2230.575 ;
        RECT 1303.720 2098.060 1304.620 2610.740 ;
        RECT 1307.020 2098.060 1371.320 2610.740 ;
        RECT 1237.020 2010.740 1371.320 2098.060 ;
        RECT 1237.020 1676.865 1301.320 2010.740 ;
        RECT 1167.020 1630.575 1301.320 1676.865 ;
        RECT 1167.020 1076.865 1231.320 1630.575 ;
        RECT 1233.720 1076.865 1234.620 1630.575 ;
        RECT 1237.020 1498.060 1301.320 1630.575 ;
        RECT 1303.720 1498.060 1304.620 2010.740 ;
        RECT 1307.020 1498.060 1371.320 2010.740 ;
        RECT 1237.020 1410.740 1371.320 1498.060 ;
        RECT 1237.020 1076.865 1301.320 1410.740 ;
        RECT 1167.020 1030.575 1301.320 1076.865 ;
        RECT 1167.020 191.935 1231.320 1030.575 ;
        RECT 1233.720 191.935 1234.620 1030.575 ;
        RECT 1237.020 898.060 1301.320 1030.575 ;
        RECT 1303.720 898.060 1304.620 1410.740 ;
        RECT 1307.020 898.060 1371.320 1410.740 ;
        RECT 1237.020 810.740 1371.320 898.060 ;
        RECT 1237.020 191.935 1301.320 810.740 ;
        RECT 1303.720 191.935 1304.620 810.740 ;
        RECT 1307.020 191.935 1371.320 810.740 ;
        RECT 1373.720 191.935 1374.620 3286.945 ;
        RECT 1377.020 2683.665 1441.320 3286.945 ;
        RECT 1443.720 2683.665 1444.620 3286.945 ;
        RECT 1447.020 2683.665 1511.320 3286.945 ;
        RECT 1377.020 2612.215 1511.320 2683.665 ;
        RECT 1377.020 2283.665 1441.320 2612.215 ;
        RECT 1443.720 2283.665 1444.620 2612.215 ;
        RECT 1447.020 2283.665 1511.320 2612.215 ;
        RECT 1377.020 2206.095 1511.320 2283.665 ;
        RECT 1377.020 2083.665 1441.320 2206.095 ;
        RECT 1443.720 2083.665 1444.620 2206.095 ;
        RECT 1447.020 2083.665 1511.320 2206.095 ;
        RECT 1377.020 2012.215 1511.320 2083.665 ;
        RECT 1377.020 1683.665 1441.320 2012.215 ;
        RECT 1443.720 1683.665 1444.620 2012.215 ;
        RECT 1447.020 1683.665 1511.320 2012.215 ;
        RECT 1377.020 1606.095 1511.320 1683.665 ;
        RECT 1377.020 1483.665 1441.320 1606.095 ;
        RECT 1443.720 1483.665 1444.620 1606.095 ;
        RECT 1447.020 1483.665 1511.320 1606.095 ;
        RECT 1377.020 1412.215 1511.320 1483.665 ;
        RECT 1377.020 1083.665 1441.320 1412.215 ;
        RECT 1443.720 1083.665 1444.620 1412.215 ;
        RECT 1447.020 1083.665 1511.320 1412.215 ;
        RECT 1377.020 1006.095 1511.320 1083.665 ;
        RECT 1377.020 883.665 1441.320 1006.095 ;
        RECT 1443.720 883.665 1444.620 1006.095 ;
        RECT 1447.020 883.665 1511.320 1006.095 ;
        RECT 1377.020 812.215 1511.320 883.665 ;
        RECT 1377.020 191.935 1441.320 812.215 ;
        RECT 1443.720 191.935 1444.620 812.215 ;
        RECT 1447.020 191.935 1511.320 812.215 ;
        RECT 1513.720 191.935 1514.620 3286.945 ;
        RECT 1517.020 191.935 1581.320 3286.945 ;
        RECT 1583.720 191.935 1584.620 3286.945 ;
        RECT 1587.020 2889.785 1651.320 3286.945 ;
        RECT 1653.720 2889.785 1654.620 3286.945 ;
        RECT 1657.020 2889.785 1721.320 3286.945 ;
        RECT 1587.020 2836.695 1721.320 2889.785 ;
        RECT 1587.020 2276.865 1651.320 2836.695 ;
        RECT 1653.720 2698.060 1654.620 2836.695 ;
        RECT 1657.020 2698.060 1721.320 2836.695 ;
        RECT 1653.720 2610.740 1721.320 2698.060 ;
        RECT 1653.720 2276.865 1654.620 2610.740 ;
        RECT 1657.020 2276.865 1721.320 2610.740 ;
        RECT 1587.020 2230.575 1721.320 2276.865 ;
        RECT 1587.020 1676.865 1651.320 2230.575 ;
        RECT 1653.720 2098.060 1654.620 2230.575 ;
        RECT 1657.020 2098.060 1721.320 2230.575 ;
        RECT 1653.720 2010.740 1721.320 2098.060 ;
        RECT 1653.720 1676.865 1654.620 2010.740 ;
        RECT 1657.020 1676.865 1721.320 2010.740 ;
        RECT 1587.020 1630.575 1721.320 1676.865 ;
        RECT 1587.020 1076.865 1651.320 1630.575 ;
        RECT 1653.720 1498.060 1654.620 1630.575 ;
        RECT 1657.020 1498.060 1721.320 1630.575 ;
        RECT 1653.720 1410.740 1721.320 1498.060 ;
        RECT 1653.720 1076.865 1654.620 1410.740 ;
        RECT 1657.020 1076.865 1721.320 1410.740 ;
        RECT 1587.020 1030.575 1721.320 1076.865 ;
        RECT 1587.020 191.935 1651.320 1030.575 ;
        RECT 1653.720 898.060 1654.620 1030.575 ;
        RECT 1657.020 898.060 1721.320 1030.575 ;
        RECT 1653.720 810.740 1721.320 898.060 ;
        RECT 1653.720 191.935 1654.620 810.740 ;
        RECT 1657.020 191.935 1721.320 810.740 ;
        RECT 1723.720 191.935 1724.620 3286.945 ;
        RECT 1727.020 191.935 1791.320 3286.945 ;
        RECT 1793.720 191.935 1794.620 3286.945 ;
        RECT 1797.020 2887.180 1861.320 3286.945 ;
        RECT 1863.720 2887.180 1864.620 3286.945 ;
        RECT 1797.020 2848.985 1864.620 2887.180 ;
        RECT 1867.020 2848.985 1915.145 3286.945 ;
        RECT 1797.020 2826.495 1915.145 2848.985 ;
        RECT 1797.020 2810.740 1864.620 2826.495 ;
        RECT 1797.020 2687.180 1861.320 2810.740 ;
        RECT 1863.720 2687.180 1864.620 2810.740 ;
        RECT 1797.020 2683.665 1864.620 2687.180 ;
        RECT 1867.020 2683.665 1915.145 2826.495 ;
        RECT 1797.020 2612.215 1915.145 2683.665 ;
        RECT 1797.020 2610.740 1864.620 2612.215 ;
        RECT 1797.020 2487.180 1861.320 2610.740 ;
        RECT 1863.720 2487.180 1864.620 2610.740 ;
        RECT 1797.020 2410.740 1864.620 2487.180 ;
        RECT 1797.020 2287.180 1861.320 2410.740 ;
        RECT 1863.720 2287.180 1864.620 2410.740 ;
        RECT 1797.020 2210.740 1864.620 2287.180 ;
        RECT 1797.020 2087.180 1861.320 2210.740 ;
        RECT 1863.720 2087.180 1864.620 2210.740 ;
        RECT 1797.020 2083.665 1864.620 2087.180 ;
        RECT 1867.020 2083.665 1915.145 2612.215 ;
        RECT 1797.020 2012.215 1915.145 2083.665 ;
        RECT 1797.020 2010.740 1864.620 2012.215 ;
        RECT 1797.020 1887.180 1861.320 2010.740 ;
        RECT 1863.720 1887.180 1864.620 2010.740 ;
        RECT 1797.020 1810.740 1864.620 1887.180 ;
        RECT 1797.020 1687.180 1861.320 1810.740 ;
        RECT 1863.720 1687.180 1864.620 1810.740 ;
        RECT 1797.020 1610.740 1864.620 1687.180 ;
        RECT 1797.020 1487.180 1861.320 1610.740 ;
        RECT 1863.720 1487.180 1864.620 1610.740 ;
        RECT 1797.020 1483.665 1864.620 1487.180 ;
        RECT 1867.020 1483.665 1915.145 2012.215 ;
        RECT 1797.020 1412.215 1915.145 1483.665 ;
        RECT 1797.020 1410.740 1864.620 1412.215 ;
        RECT 1797.020 1287.180 1861.320 1410.740 ;
        RECT 1863.720 1287.180 1864.620 1410.740 ;
        RECT 1797.020 1210.740 1864.620 1287.180 ;
        RECT 1797.020 1087.180 1861.320 1210.740 ;
        RECT 1863.720 1087.180 1864.620 1210.740 ;
        RECT 1797.020 1010.740 1864.620 1087.180 ;
        RECT 1797.020 887.180 1861.320 1010.740 ;
        RECT 1863.720 887.180 1864.620 1010.740 ;
        RECT 1797.020 883.665 1864.620 887.180 ;
        RECT 1867.020 883.665 1915.145 1412.215 ;
        RECT 1797.020 812.215 1915.145 883.665 ;
        RECT 1797.020 810.740 1864.620 812.215 ;
        RECT 1797.020 687.180 1861.320 810.740 ;
        RECT 1863.720 687.180 1864.620 810.740 ;
        RECT 1797.020 610.740 1864.620 687.180 ;
        RECT 1797.020 487.180 1861.320 610.740 ;
        RECT 1863.720 487.180 1864.620 610.740 ;
        RECT 1797.020 410.740 1864.620 487.180 ;
        RECT 1797.020 191.935 1861.320 410.740 ;
        RECT 1863.720 191.935 1864.620 410.740 ;
        RECT 1867.020 191.935 1915.145 812.215 ;
  END
END user_proj_example
END LIBRARY

